
module biquad_filter ( clk, en, reset, \parameter_A1_mul[7] , 
        \parameter_A1_mul[6] , \parameter_A1_mul[5] , \parameter_A1_mul[4] , 
        \parameter_A1_mul[3] , \parameter_A1_mul[2] , \parameter_A1_mul[1] , 
        \parameter_A1_mul[0] , \parameter_A1_div[7] , \parameter_A1_div[6] , 
        \parameter_A1_div[5] , \parameter_A1_div[4] , \parameter_A1_div[3] , 
        \parameter_A1_div[2] , \parameter_A1_div[1] , \parameter_A1_div[0] , 
        \parameter_A2_mul[7] , \parameter_A2_mul[6] , \parameter_A2_mul[5] , 
        \parameter_A2_mul[4] , \parameter_A2_mul[3] , \parameter_A2_mul[2] , 
        \parameter_A2_mul[1] , \parameter_A2_mul[0] , \parameter_A2_div[7] , 
        \parameter_A2_div[6] , \parameter_A2_div[5] , \parameter_A2_div[4] , 
        \parameter_A2_div[3] , \parameter_A2_div[2] , \parameter_A2_div[1] , 
        \parameter_A2_div[0] , \parameter_B0_mul[7] , \parameter_B0_mul[6] , 
        \parameter_B0_mul[5] , \parameter_B0_mul[4] , \parameter_B0_mul[3] , 
        \parameter_B0_mul[2] , \parameter_B0_mul[1] , \parameter_B0_mul[0] , 
        \parameter_B0_div[7] , \parameter_B0_div[6] , \parameter_B0_div[5] , 
        \parameter_B0_div[4] , \parameter_B0_div[3] , \parameter_B0_div[2] , 
        \parameter_B0_div[1] , \parameter_B0_div[0] , \parameter_B1_mul[7] , 
        \parameter_B1_mul[6] , \parameter_B1_mul[5] , \parameter_B1_mul[4] , 
        \parameter_B1_mul[3] , \parameter_B1_mul[2] , \parameter_B1_mul[1] , 
        \parameter_B1_mul[0] , \parameter_B1_div[7] , \parameter_B1_div[6] , 
        \parameter_B1_div[5] , \parameter_B1_div[4] , \parameter_B1_div[3] , 
        \parameter_B1_div[2] , \parameter_B1_div[1] , \parameter_B1_div[0] , 
        \parameter_B2_mul[7] , \parameter_B2_mul[6] , \parameter_B2_mul[5] , 
        \parameter_B2_mul[4] , \parameter_B2_mul[3] , \parameter_B2_mul[2] , 
        \parameter_B2_mul[1] , \parameter_B2_mul[0] , \parameter_B2_div[7] , 
        \parameter_B2_div[6] , \parameter_B2_div[5] , \parameter_B2_div[4] , 
        \parameter_B2_div[3] , \parameter_B2_div[2] , \parameter_B2_div[1] , 
        \parameter_B2_div[0] , \input_signal[7] , \input_signal[6] , 
        \input_signal[5] , \input_signal[4] , \input_signal[3] , 
        \input_signal[2] , \input_signal[1] , \input_signal[0] , 
        \output_signal[7] , \output_signal[6] , \output_signal[5] , 
        \output_signal[4] , \output_signal[3] , \output_signal[2] , 
        \output_signal[1] , \output_signal[0] , change_input, 
        temporary_overflow );
  input clk, en, reset, \parameter_A1_mul[7] , \parameter_A1_mul[6] ,
         \parameter_A1_mul[5] , \parameter_A1_mul[4] , \parameter_A1_mul[3] ,
         \parameter_A1_mul[2] , \parameter_A1_mul[1] , \parameter_A1_mul[0] ,
         \parameter_A1_div[7] , \parameter_A1_div[6] , \parameter_A1_div[5] ,
         \parameter_A1_div[4] , \parameter_A1_div[3] , \parameter_A1_div[2] ,
         \parameter_A1_div[1] , \parameter_A1_div[0] , \parameter_A2_mul[7] ,
         \parameter_A2_mul[6] , \parameter_A2_mul[5] , \parameter_A2_mul[4] ,
         \parameter_A2_mul[3] , \parameter_A2_mul[2] , \parameter_A2_mul[1] ,
         \parameter_A2_mul[0] , \parameter_A2_div[7] , \parameter_A2_div[6] ,
         \parameter_A2_div[5] , \parameter_A2_div[4] , \parameter_A2_div[3] ,
         \parameter_A2_div[2] , \parameter_A2_div[1] , \parameter_A2_div[0] ,
         \parameter_B0_mul[7] , \parameter_B0_mul[6] , \parameter_B0_mul[5] ,
         \parameter_B0_mul[4] , \parameter_B0_mul[3] , \parameter_B0_mul[2] ,
         \parameter_B0_mul[1] , \parameter_B0_mul[0] , \parameter_B0_div[7] ,
         \parameter_B0_div[6] , \parameter_B0_div[5] , \parameter_B0_div[4] ,
         \parameter_B0_div[3] , \parameter_B0_div[2] , \parameter_B0_div[1] ,
         \parameter_B0_div[0] , \parameter_B1_mul[7] , \parameter_B1_mul[6] ,
         \parameter_B1_mul[5] , \parameter_B1_mul[4] , \parameter_B1_mul[3] ,
         \parameter_B1_mul[2] , \parameter_B1_mul[1] , \parameter_B1_mul[0] ,
         \parameter_B1_div[7] , \parameter_B1_div[6] , \parameter_B1_div[5] ,
         \parameter_B1_div[4] , \parameter_B1_div[3] , \parameter_B1_div[2] ,
         \parameter_B1_div[1] , \parameter_B1_div[0] , \parameter_B2_mul[7] ,
         \parameter_B2_mul[6] , \parameter_B2_mul[5] , \parameter_B2_mul[4] ,
         \parameter_B2_mul[3] , \parameter_B2_mul[2] , \parameter_B2_mul[1] ,
         \parameter_B2_mul[0] , \parameter_B2_div[7] , \parameter_B2_div[6] ,
         \parameter_B2_div[5] , \parameter_B2_div[4] , \parameter_B2_div[3] ,
         \parameter_B2_div[2] , \parameter_B2_div[1] , \parameter_B2_div[0] ,
         \input_signal[7] , \input_signal[6] , \input_signal[5] ,
         \input_signal[4] , \input_signal[3] , \input_signal[2] ,
         \input_signal[1] , \input_signal[0] ;
  output \output_signal[7] , \output_signal[6] , \output_signal[5] ,
         \output_signal[4] , \output_signal[3] , \output_signal[2] ,
         \output_signal[1] , \output_signal[0] , change_input,
         temporary_overflow;
  wire   n4673, output_contracterxn8, output_contracterxn7,
         output_contracterxn6, output_contracterxn5, output_contracterxn4,
         output_contracterxn3, output_contracterxn2, output_contracterxn1,
         input_prev_0_registerxn20, input_prev_0_registerxn18,
         input_prev_0_registerxn17, input_prev_0_registerxn16,
         input_prev_0_registerxn15, input_prev_0_registerxn14,
         input_prev_0_registerxn13, input_prev_0_registerxn12,
         input_prev_0_registerxn11, input_prev_0_registerxn10,
         input_prev_0_registerxn9, input_prev_0_registerxn8,
         input_prev_0_registerxn7, input_prev_0_registerxn6,
         input_prev_0_registerxn5, input_prev_0_registerxn4,
         input_prev_0_registerxn3, input_prev_0_registerxn2,
         input_times_b0_mul_componentxn108, input_times_b0_mul_componentxn107,
         input_times_b0_mul_componentxn106, input_times_b0_mul_componentxn105,
         input_times_b0_mul_componentxn104, input_times_b0_mul_componentxn103,
         input_times_b0_mul_componentxn102, input_times_b0_mul_componentxn101,
         input_times_b0_mul_componentxn100, input_times_b0_mul_componentxn99,
         input_times_b0_mul_componentxn98, input_times_b0_mul_componentxn97,
         input_times_b0_mul_componentxn96, input_times_b0_mul_componentxn95,
         input_times_b0_mul_componentxn94, input_times_b0_mul_componentxn93,
         input_times_b0_mul_componentxn92, input_times_b0_mul_componentxn91,
         input_times_b0_mul_componentxn90, input_times_b0_mul_componentxn89,
         input_times_b0_mul_componentxn88, input_times_b0_mul_componentxn87,
         input_times_b0_mul_componentxn86, input_times_b0_mul_componentxn85,
         input_times_b0_mul_componentxn84, input_times_b0_mul_componentxn83,
         input_times_b0_mul_componentxn82, input_times_b0_mul_componentxn81,
         input_times_b0_mul_componentxn80, input_times_b0_mul_componentxn79,
         input_times_b0_mul_componentxn78, input_times_b0_mul_componentxn77,
         input_times_b0_mul_componentxn76, input_times_b0_mul_componentxn75,
         input_times_b0_mul_componentxn74, input_times_b0_mul_componentxn73,
         input_times_b0_mul_componentxn72, input_times_b0_mul_componentxn71,
         input_times_b0_mul_componentxn70, input_times_b0_mul_componentxn69,
         input_times_b0_mul_componentxn68, input_times_b0_mul_componentxn67,
         input_times_b0_mul_componentxn66, input_times_b0_mul_componentxn65,
         input_times_b0_mul_componentxn64, input_times_b0_mul_componentxn63,
         input_times_b0_mul_componentxn62, input_times_b0_mul_componentxn61,
         input_times_b0_mul_componentxn60, input_times_b0_mul_componentxn59,
         input_times_b0_mul_componentxn58, input_times_b0_mul_componentxn57,
         input_times_b0_mul_componentxn56,
         input_times_b0_mul_componentxunsigned_output_8,
         input_times_b0_mul_componentxunsigned_output_9,
         input_times_b0_mul_componentxunsigned_output_10,
         input_times_b0_mul_componentxunsigned_output_11,
         input_times_b0_mul_componentxunsigned_output_12,
         input_times_b0_mul_componentxunsigned_output_13,
         input_times_b0_mul_componentxunsigned_output_14,
         input_times_b0_mul_componentxunsigned_output_15,
         input_times_b0_mul_componentxunsigned_output_16,
         input_times_b0_mul_componentxunsigned_output_17,
         input_times_b0_mul_componentxinput_B_inverted_1_,
         input_times_b0_mul_componentxinput_B_inverted_2_,
         input_times_b0_mul_componentxinput_B_inverted_3_,
         input_times_b0_mul_componentxinput_B_inverted_4_,
         input_times_b0_mul_componentxinput_B_inverted_5_,
         input_times_b0_mul_componentxinput_B_inverted_6_,
         input_times_b0_mul_componentxinput_B_inverted_7_,
         input_times_b0_mul_componentxinput_B_inverted_8_,
         input_times_b0_mul_componentxinput_B_inverted_9_,
         input_times_b0_mul_componentxinput_B_inverted_10_,
         input_times_b0_mul_componentxinput_B_inverted_11_,
         input_times_b0_mul_componentxinput_B_inverted_12_,
         input_times_b0_mul_componentxinput_B_inverted_13_,
         input_times_b0_mul_componentxinput_B_inverted_14_,
         input_times_b0_mul_componentxinput_B_inverted_15_,
         input_times_b0_mul_componentxinput_B_inverted_16_,
         input_times_b0_mul_componentxinput_B_inverted_17_,
         input_times_b0_div_componentxn62, input_times_b0_div_componentxn61,
         input_times_b0_div_componentxn60, input_times_b0_div_componentxn59,
         input_times_b0_div_componentxn58, input_times_b0_div_componentxn57,
         input_times_b0_div_componentxn56, input_times_b0_div_componentxn55,
         input_times_b0_div_componentxn54, input_times_b0_div_componentxn53,
         input_times_b0_div_componentxn52, input_times_b0_div_componentxn51,
         input_times_b0_div_componentxn50, input_times_b0_div_componentxn49,
         input_times_b0_div_componentxn48, input_times_b0_div_componentxn47,
         input_times_b0_div_componentxn46, input_times_b0_div_componentxn45,
         input_times_b0_div_componentxn44, input_times_b0_div_componentxn43,
         input_times_b0_div_componentxn42, input_times_b0_div_componentxn41,
         input_times_b0_div_componentxn40, input_times_b0_div_componentxn39,
         input_times_b0_div_componentxn38, input_times_b0_div_componentxn37,
         input_times_b0_div_componentxn36, input_times_b0_div_componentxn35,
         input_times_b0_div_componentxn34, input_times_b0_div_componentxn33,
         input_times_b0_div_componentxn32, input_times_b0_div_componentxn31,
         input_times_b0_div_componentxn30, input_times_b0_div_componentxn29,
         input_times_b0_div_componentxn28, input_times_b0_div_componentxn27,
         input_times_b0_div_componentxn25, input_times_b0_div_componentxn24,
         input_times_b0_div_componentxn21, input_times_b0_div_componentxn20,
         input_times_b0_div_componentxn19, input_times_b0_div_componentxn18,
         input_times_b0_div_componentxn17, input_times_b0_div_componentxn16,
         input_times_b0_div_componentxn15, input_times_b0_div_componentxn14,
         input_times_b0_div_componentxn13, input_times_b0_div_componentxn12,
         input_times_b0_div_componentxn11, input_times_b0_div_componentxn10,
         input_times_b0_div_componentxn9, input_times_b0_div_componentxn8,
         input_times_b0_div_componentxn7, input_times_b0_div_componentxn6,
         input_times_b0_div_componentxn5, input_times_b0_div_componentxn3,
         input_times_b0_div_componentxoutput_sign_gated,
         input_times_b0_div_componentxoutput_sign_gated_prev,
         input_times_b0_div_componentxunsigned_B_17,
         input_times_b0_div_componentxunsigned_A_17,
         input_times_b0_div_componentxunsigned_output_1,
         input_times_b0_div_componentxunsigned_output_2,
         input_times_b0_div_componentxunsigned_output_3,
         input_times_b0_div_componentxunsigned_output_4,
         input_times_b0_div_componentxunsigned_output_5,
         input_times_b0_div_componentxunsigned_output_6,
         input_times_b0_div_componentxunsigned_output_7,
         input_times_b0_div_componentxunsigned_output_8,
         input_times_b0_div_componentxunsigned_output_9,
         input_times_b0_div_componentxunsigned_output_10,
         input_times_b0_div_componentxunsigned_output_11,
         input_times_b0_div_componentxunsigned_output_12,
         input_times_b0_div_componentxunsigned_output_13,
         input_times_b0_div_componentxunsigned_output_14,
         input_times_b0_div_componentxunsigned_output_15,
         input_times_b0_div_componentxunsigned_output_16,
         input_times_b0_div_componentxunsigned_output_17,
         input_times_b0_div_componentxinput_B_inverted_1_,
         input_times_b0_div_componentxinput_B_inverted_2_,
         input_times_b0_div_componentxinput_B_inverted_3_,
         input_times_b0_div_componentxinput_B_inverted_4_,
         input_times_b0_div_componentxinput_B_inverted_5_,
         input_times_b0_div_componentxinput_B_inverted_6_,
         input_times_b0_div_componentxinput_B_inverted_7_,
         input_times_b0_div_componentxinput_B_inverted_8_,
         input_times_b0_div_componentxinput_B_inverted_9_,
         input_times_b0_div_componentxinput_B_inverted_10_,
         input_times_b0_div_componentxinput_B_inverted_11_,
         input_times_b0_div_componentxinput_B_inverted_12_,
         input_times_b0_div_componentxinput_B_inverted_13_,
         input_times_b0_div_componentxinput_B_inverted_14_,
         input_times_b0_div_componentxinput_B_inverted_15_,
         input_times_b0_div_componentxinput_B_inverted_16_,
         input_times_b0_div_componentxinput_B_inverted_17_,
         results_b0_b1_adderxn35, results_b0_b1_adderxn34,
         results_b0_b1_adderxn33, results_b0_b1_adderxn32,
         results_b0_b1_adderxn31, results_b0_b1_adderxn30,
         results_b0_b1_adderxn29, results_b0_b1_adderxn28,
         results_b0_b1_adderxn27, results_b0_b1_adderxn26,
         results_b0_b1_adderxn25, results_b0_b1_adderxn24,
         results_b0_b1_adderxn23, results_b0_b1_adderxn22,
         results_b0_b1_adderxn21, results_b0_b1_adderxn20,
         results_b0_b1_adderxn19, results_b0_b1_adderxn17,
         results_b0_b1_adderxn16, results_b0_b1_adderxn15,
         results_b0_b1_adderxn14, results_b0_b1_adderxn13,
         results_b0_b1_adderxn12, results_b0_b1_adderxn11,
         results_b0_b1_adderxn10, results_b0_b1_adderxn9,
         results_b0_b1_adderxn8, results_b0_b1_adderxn7,
         results_b0_b1_adderxn6, results_b0_b1_adderxn5,
         results_b0_b1_adderxn4, results_b0_b1_adderxn3,
         results_b0_b1_adderxn2, results_a1_a2_inv_inverterxn17,
         results_a1_a2_inv_inverterxn15, results_a1_a2_inv_inverterxn13,
         results_a1_a2_inv_inverterxn12, results_a1_a2_inv_inverterxn11,
         results_a1_a2_inv_inverterxn10, results_a1_a2_inv_inverterxn9,
         results_a1_a2_inv_inverterxn8, results_a1_a2_inv_inverterxn6,
         results_a1_a2_inv_inverterxn4, results_a1_a2_inv_inverterxn2,
         clock_chopper_and_divisionxn49, clock_chopper_and_divisionxn47,
         clock_chopper_and_divisionxn46, clock_chopper_and_divisionxn45,
         clock_chopper_and_divisionxn44, clock_chopper_and_divisionxn43,
         clock_chopper_and_divisionxn42, clock_chopper_and_divisionxn41,
         clock_chopper_and_divisionxn40, clock_chopper_and_divisionxn39,
         clock_chopper_and_divisionxn38, clock_chopper_and_divisionxn37,
         clock_chopper_and_divisionxn36, clock_chopper_and_divisionxn35,
         clock_chopper_and_divisionxn34, clock_chopper_and_divisionxn33,
         clock_chopper_and_divisionxn32, clock_chopper_and_divisionxn31,
         clock_chopper_and_divisionxn30, clock_chopper_and_divisionxn29,
         clock_chopper_and_divisionxn28, clock_chopper_and_divisionxn27,
         clock_chopper_and_divisionxn26,
         input_times_b0_mul_componentxUMxsum_layer5_128315744_128315968_128316136,
         input_times_b0_mul_componentxUMxsum_layer5_128315464_128315632_128315800,
         input_times_b0_mul_componentxUMxsum_layer5_128220800_128221024_128221136,
         input_times_b0_mul_componentxUMxsum_layer5_128220688_128220856_128220968,
         input_times_b0_mul_componentxUMxsum_layer5_128126256_128220520_128220744,
         input_times_b0_mul_componentxUMxsum_layer5_128125920_128220352_128220576,
         input_times_b0_mul_componentxUMxsum_layer5_128125584_128220184_128220408,
         input_times_b0_mul_componentxUMxsum_layer5_128125248_128219960_128220240,
         input_times_b0_mul_componentxUMxcarry_layer5_128219792_128220016,
         input_times_b0_mul_componentxUMxsum_layer5_128219792_128220016,
         input_times_b0_mul_componentxUMxcarry_layer5_128219624_128219848,
         input_times_b0_mul_componentxUMxsum_layer5_128219624_128219848,
         input_times_b0_mul_componentxUMxcarry_layer5_128219456_128219680,
         input_times_b0_mul_componentxUMxsum_layer5_128219456_128219680,
         input_times_b0_mul_componentxUMxcarry_layer5_128219288_128219512,
         input_times_b0_mul_componentxUMxsum_layer5_128219288_128219512,
         input_times_b0_mul_componentxUMxcarry_layer5_128219120_128219344,
         input_times_b0_mul_componentxUMxsum_layer4_128238312_128238424_128238592,
         input_times_b0_mul_componentxUMxsum_layer4_128237752_128237976_128238144,
         input_times_b0_mul_componentxUMxsum_layer4_128237920_128238088,
         input_times_b0_mul_componentxUMxsum_layer4_128126760_128237640_128237808,
         input_times_b0_mul_componentxUMxcarry_layer4_128126816_128126928,
         input_times_b0_mul_componentxUMxsum_layer4_128126816_128126928,
         input_times_b0_mul_componentxUMxsum_layer4_128263168_128126424_128126648,
         input_times_b0_mul_componentxUMxcarry_layer4_128126480_128126592,
         input_times_b0_mul_componentxUMxsum_layer4_128126480_128126592,
         input_times_b0_mul_componentxUMxsum_layer4_128262496_128126088_128126312,
         input_times_b0_mul_componentxUMxsum_layer4_128125752_128125976_128126144,
         input_times_b0_mul_componentxUMxsum_layer4_128125416_128125640_128125808,
         input_times_b0_mul_componentxUMxsum_layer4_128125080_128125304_128125472,
         input_times_b0_mul_componentxUMxsum_layer4_128124744_128124968_128125136,
         input_times_b0_mul_componentxUMxsum_layer4_128124632_128124800_128124912,
         input_times_b0_mul_componentxUMxsum_layer4_128247456_128124464_128124688,
         input_times_b0_mul_componentxUMxsum_layer4_128247120_128124240_128124520,
         input_times_b0_mul_componentxUMxcarry_layer4_128124072_128124296,
         input_times_b0_mul_componentxUMxsum_layer4_128124072_128124296,
         input_times_b0_mul_componentxUMxcarry_layer4_128123904_128124128,
         input_times_b0_mul_componentxUMxsum_layer4_128123904_128124128,
         input_times_b0_mul_componentxUMxcarry_layer4_128123792_128123960,
         input_times_b0_mul_componentxUMxsum_layer3_128264344_128264512,
         input_times_b0_mul_componentxUMxsum_layer3_128263896_128264064_128264176,
         input_times_b0_mul_componentxUMxsum_layer3_128263336_128263560_128263728,
         input_times_b0_mul_componentxUMxcarry_layer3_128263672_128263840,
         input_times_b0_mul_componentxUMxsum_layer3_128263672_128263840,
         input_times_b0_mul_componentxUMxsum_layer3_128263224_128263392_128263504,
         input_times_b0_mul_componentxUMxsum_layer3_128262664_128262888_128263056,
         input_times_b0_mul_componentxUMxsum_layer3_128262720_128262832_128263000,
         input_times_b0_mul_componentxUMxsum_layer3_128262216_128262384_128262552,
         input_times_b0_mul_componentxUMxsum_layer3_128249696_128249808_128262328,
         input_times_b0_mul_componentxUMxsum_layer3_128197128_128249304_128249528,
         input_times_b0_mul_componentxUMxsum_layer3_128249360_128249472_128249640,
         input_times_b0_mul_componentxUMxsum_layer3_128248800_128249024_128249192,
         input_times_b0_mul_componentxUMxsum_layer3_128248856_128248968_128249136,
         input_times_b0_mul_componentxUMxsum_layer3_128248296_128248520_128248688,
         input_times_b0_mul_componentxUMxcarry_layer3_128248464_128248632,
         input_times_b0_mul_componentxUMxsum_layer3_128248464_128248632,
         input_times_b0_mul_componentxUMxsum_layer3_128247960_128248184_128248352,
         input_times_b0_mul_componentxUMxcarry_layer3_128248016_128248128,
         input_times_b0_mul_componentxUMxsum_layer3_128248016_128248128,
         input_times_b0_mul_componentxUMxsum_layer3_128222880_128247624_128247848,
         input_times_b0_mul_componentxUMxcarry_layer3_128247680_128247792,
         input_times_b0_mul_componentxUMxsum_layer3_128247680_128247792,
         input_times_b0_mul_componentxUMxsum_layer3_128222208_128247288_128247512,
         input_times_b0_mul_componentxUMxsum_layer3_128246952_128247176_128247344,
         input_times_b0_mul_componentxUMxsum_layer3_128246616_128246840_128247008,
         input_times_b0_mul_componentxUMxsum_layer3_128246504_128246672_128246784,
         input_times_b0_mul_componentxUMxsum_layer3_127827080_128246280_128246560,
         input_times_b0_mul_componentxUMxcarry_layer3_128246112_128246336,
         input_times_b0_mul_componentxUMxsum_layer3_128246112_128246336,
         input_times_b0_mul_componentxUMxcarry_layer3_128246000_128246168,
         input_times_b0_mul_componentxUMxsum_layer2_128199816_128200040_128199984,
         input_times_b0_mul_componentxUMxsum_layer2_128199368_128199480_128199648,
         input_times_b0_mul_componentxUMxsum_layer2_128198864_128199032_128199200,
         input_times_b0_mul_componentxUMxsum_layer2_128198304_128198528_128198696,
         input_times_b0_mul_componentxUMxcarry_layer2_128198976_128199144,
         input_times_b0_mul_componentxUMxsum_layer2_128198976_128199144,
         input_times_b0_mul_componentxUMxsum_layer2_128198472_128198640_128198808,
         input_times_b0_mul_componentxUMxsum_layer2_128198080_128198192_128198360,
         input_times_b0_mul_componentxUMxsum_layer2_128197464_128197688_128197856,
         input_times_b0_mul_componentxUMxcarry_layer2_128198024_128197968,
         input_times_b0_mul_componentxUMxsum_layer2_128198024_128197968,
         input_times_b0_mul_componentxUMxsum_layer2_128197520_128197632_128197800,
         input_times_b0_mul_componentxUMxsum_layer2_128197016_128197240_128197352,
         input_times_b0_mul_componentxUMxsum_layer2_127627392_128196680_128196848,
         input_times_b0_mul_componentxUMxa15_and_b0,
         input_times_b0_mul_componentxUMxsum_layer2_128196792_128196960_128197184,
         input_times_b0_mul_componentxUMxsum_layer2_128224952_128225120_128225232,
         input_times_b0_mul_componentxUMxsum_layer2_128224392_128224616_128224784,
         input_times_b0_mul_componentxUMxsum_layer2_128224728_128224896_128225064,
         input_times_b0_mul_componentxUMxsum_layer2_128224280_128224448_128224560,
         input_times_b0_mul_componentxUMxsum_layer2_128223720_128223944_128224168,
         input_times_b0_mul_componentxUMxsum_layer2_128223888_128224112_128224056,
         input_times_b0_mul_componentxUMxsum_layer2_128223440_128223608_128223776,
         input_times_b0_mul_componentxUMxsum_layer2_127715424_128223048_128223272,
         input_times_b0_mul_componentxUMxa12_and_b0,
         input_times_b0_mul_componentxUMxcarry_layer2_128223384_128223552,
         input_times_b0_mul_componentxUMxsum_layer2_128223384_128223552,
         input_times_b0_mul_componentxUMxsum_layer2_128222936_128223104_128223216,
         input_times_b0_mul_componentxUMxsum_layer2_128222376_128222600_128222768,
         input_times_b0_mul_componentxUMxsum_layer2_128222432_128222544_128222712,
         input_times_b0_mul_componentxUMxsum_layer2_128221872_128222096_128222264,
         input_times_b0_mul_componentxUMxsum_layer2_128221760_128221928_128222040,
         input_times_b0_mul_componentxUMxsum_layer2_127635584_128221368_128221592,
         input_times_b0_mul_componentxUMxa9_and_b0,
         input_times_b0_mul_componentxUMxsum_layer2_128221424_128221536_128221704,
         input_times_b0_mul_componentxUMxsum_layer2_127827584_127827808_128221256,
         input_times_b0_mul_componentxUMxcarry_layer2_127827752_127827920,
         input_times_b0_mul_componentxUMxsum_layer2_127827752_127827920,
         input_times_b0_mul_componentxUMxsum_layer2_127827248_127827472_127827640,
         input_times_b0_mul_componentxUMxcarry_layer2_127827304_127827416,
         input_times_b0_mul_componentxUMxsum_layer2_127827304_127827416,
         input_times_b0_mul_componentxUMxsum_layer2_127731808_127826912_127827136,
         input_times_b0_mul_componentxUMxa6_and_b0,
         input_times_b0_mul_componentxUMxsum_layer2_127826576_127826800_127826968,
         input_times_b0_mul_componentxUMxsum_layer2_127826464_127826632_127826744,
         input_times_b0_mul_componentxUMxsum_layer2_127672448_127826240_127826520,
         input_times_b0_mul_componentxUMxa3_and_b0,
         input_times_b0_mul_componentxUMxcarry_layer2_127826128_127826296,
         input_times_b0_mul_componentxUMxsum_layer1_127627616_127629520_127824000,
         input_times_b0_mul_componentxUMxa17_and_b0,
         input_times_b0_mul_componentxUMxa16_and_b1,
         input_times_b0_mul_componentxUMxa15_and_b2,
         input_times_b0_mul_componentxUMxsum_layer1_127715984_127849024_127850928,
         input_times_b0_mul_componentxUMxa14_and_b3,
         input_times_b0_mul_componentxUMxa13_and_b4,
         input_times_b0_mul_componentxUMxa12_and_b5,
         input_times_b0_mul_componentxUMxsum_layer1_127636480_127638384_127714080,
         input_times_b0_mul_componentxUMxa11_and_b6,
         input_times_b0_mul_componentxUMxa10_and_b7,
         input_times_b0_mul_componentxUMxa9_and_b8,
         input_times_b0_mul_componentxUMxsum_layer1_127733040_127722720_127724624,
         input_times_b0_mul_componentxUMxa8_and_b9,
         input_times_b0_mul_componentxUMxa7_and_b10,
         input_times_b0_mul_componentxUMxa6_and_b11,
         input_times_b0_mul_componentxUMxsum_layer1_127674016_127675920_127731136,
         input_times_b0_mul_componentxUMxa5_and_b12,
         input_times_b0_mul_componentxUMxa4_and_b13,
         input_times_b0_mul_componentxUMxa3_and_b14,
         input_times_b0_mul_componentxUMxsum_layer1_127832016_127846272_127848176,
         input_times_b0_mul_componentxUMxa2_and_b15,
         input_times_b0_mul_componentxUMxa1_and_b16,
         input_times_b0_mul_componentxUMxa0_and_b17,
         input_times_b0_mul_componentxUMxcarry_layer1_127627504_127629408,
         input_times_b0_mul_componentxUMxsum_layer1_127627504_127629408,
         input_times_b0_mul_componentxUMxa16_and_b0,
         input_times_b0_mul_componentxUMxa15_and_b1,
         input_times_b0_mul_componentxUMxsum_layer1_127715872_127848912_127850816,
         input_times_b0_mul_componentxUMxa14_and_b2,
         input_times_b0_mul_componentxUMxa13_and_b3,
         input_times_b0_mul_componentxUMxa12_and_b4,
         input_times_b0_mul_componentxUMxsum_layer1_127636368_127638272_127713968,
         input_times_b0_mul_componentxUMxa11_and_b5,
         input_times_b0_mul_componentxUMxa10_and_b6,
         input_times_b0_mul_componentxUMxa9_and_b7,
         input_times_b0_mul_componentxUMxsum_layer1_127732928_127722608_127724512,
         input_times_b0_mul_componentxUMxa8_and_b8,
         input_times_b0_mul_componentxUMxa7_and_b9,
         input_times_b0_mul_componentxUMxa6_and_b10,
         input_times_b0_mul_componentxUMxsum_layer1_127673904_127675808_127731024,
         input_times_b0_mul_componentxUMxa5_and_b11,
         input_times_b0_mul_componentxUMxa4_and_b12,
         input_times_b0_mul_componentxUMxa3_and_b13,
         input_times_b0_mul_componentxUMxsum_layer1_127831904_127846160_127848064,
         input_times_b0_mul_componentxUMxa2_and_b14,
         input_times_b0_mul_componentxUMxa1_and_b15,
         input_times_b0_mul_componentxUMxa0_and_b16,
         input_times_b0_mul_componentxUMxsum_layer1_127715760_127848800_127850704,
         input_times_b0_mul_componentxUMxa14_and_b1,
         input_times_b0_mul_componentxUMxa13_and_b2,
         input_times_b0_mul_componentxUMxa12_and_b3,
         input_times_b0_mul_componentxUMxsum_layer1_127636256_127638160_127713856,
         input_times_b0_mul_componentxUMxa11_and_b4,
         input_times_b0_mul_componentxUMxa10_and_b5,
         input_times_b0_mul_componentxUMxa9_and_b6,
         input_times_b0_mul_componentxUMxsum_layer1_127732816_127722496_127724400,
         input_times_b0_mul_componentxUMxa8_and_b7,
         input_times_b0_mul_componentxUMxa7_and_b8,
         input_times_b0_mul_componentxUMxa6_and_b9,
         input_times_b0_mul_componentxUMxsum_layer1_127673792_127675696_127730912,
         input_times_b0_mul_componentxUMxa5_and_b10,
         input_times_b0_mul_componentxUMxa4_and_b11,
         input_times_b0_mul_componentxUMxa3_and_b12,
         input_times_b0_mul_componentxUMxsum_layer1_127831792_127846048_127847952,
         input_times_b0_mul_componentxUMxa2_and_b13,
         input_times_b0_mul_componentxUMxa1_and_b14,
         input_times_b0_mul_componentxUMxa0_and_b15,
         input_times_b0_mul_componentxUMxsum_layer1_127715648_127848688_127850592,
         input_times_b0_mul_componentxUMxa14_and_b0,
         input_times_b0_mul_componentxUMxa13_and_b1,
         input_times_b0_mul_componentxUMxa12_and_b2,
         input_times_b0_mul_componentxUMxsum_layer1_127636144_127638048_127713744,
         input_times_b0_mul_componentxUMxa11_and_b3,
         input_times_b0_mul_componentxUMxa10_and_b4,
         input_times_b0_mul_componentxUMxa9_and_b5,
         input_times_b0_mul_componentxUMxsum_layer1_127732704_127722384_127724288,
         input_times_b0_mul_componentxUMxa8_and_b6,
         input_times_b0_mul_componentxUMxa7_and_b7,
         input_times_b0_mul_componentxUMxa6_and_b8,
         input_times_b0_mul_componentxUMxsum_layer1_127673680_127675584_127730800,
         input_times_b0_mul_componentxUMxa5_and_b9,
         input_times_b0_mul_componentxUMxa4_and_b10,
         input_times_b0_mul_componentxUMxa3_and_b11,
         input_times_b0_mul_componentxUMxsum_layer1_127831680_127845936_127847840,
         input_times_b0_mul_componentxUMxa2_and_b12,
         input_times_b0_mul_componentxUMxa1_and_b13,
         input_times_b0_mul_componentxUMxa0_and_b14,
         input_times_b0_mul_componentxUMxcarry_layer1_127715536_127848576,
         input_times_b0_mul_componentxUMxsum_layer1_127715536_127848576,
         input_times_b0_mul_componentxUMxa13_and_b0,
         input_times_b0_mul_componentxUMxa12_and_b1,
         input_times_b0_mul_componentxUMxsum_layer1_127636032_127637936_127713632,
         input_times_b0_mul_componentxUMxa11_and_b2,
         input_times_b0_mul_componentxUMxa10_and_b3,
         input_times_b0_mul_componentxUMxa9_and_b4,
         input_times_b0_mul_componentxUMxsum_layer1_127732592_127722272_127724176,
         input_times_b0_mul_componentxUMxa8_and_b5,
         input_times_b0_mul_componentxUMxa7_and_b6,
         input_times_b0_mul_componentxUMxa6_and_b7,
         input_times_b0_mul_componentxUMxsum_layer1_127673568_127675472_127730688,
         input_times_b0_mul_componentxUMxa5_and_b8,
         input_times_b0_mul_componentxUMxa4_and_b9,
         input_times_b0_mul_componentxUMxa3_and_b10,
         input_times_b0_mul_componentxUMxsum_layer1_127831568_127845824_127847728,
         input_times_b0_mul_componentxUMxa2_and_b11,
         input_times_b0_mul_componentxUMxa1_and_b12,
         input_times_b0_mul_componentxUMxa0_and_b13,
         input_times_b0_mul_componentxUMxsum_layer1_127635920_127637824_127713520,
         input_times_b0_mul_componentxUMxa11_and_b1,
         input_times_b0_mul_componentxUMxa10_and_b2,
         input_times_b0_mul_componentxUMxa9_and_b3,
         input_times_b0_mul_componentxUMxsum_layer1_127732480_127722160_127724064,
         input_times_b0_mul_componentxUMxa8_and_b4,
         input_times_b0_mul_componentxUMxa7_and_b5,
         input_times_b0_mul_componentxUMxa6_and_b6,
         input_times_b0_mul_componentxUMxsum_layer1_127673456_127675360_127730576,
         input_times_b0_mul_componentxUMxa5_and_b7,
         input_times_b0_mul_componentxUMxa4_and_b8,
         input_times_b0_mul_componentxUMxa3_and_b9,
         input_times_b0_mul_componentxUMxsum_layer1_127831456_127845712_127847616,
         input_times_b0_mul_componentxUMxa2_and_b10,
         input_times_b0_mul_componentxUMxa1_and_b11,
         input_times_b0_mul_componentxUMxa0_and_b12,
         input_times_b0_mul_componentxUMxsum_layer1_127635808_127637712_127713408,
         input_times_b0_mul_componentxUMxa11_and_b0,
         input_times_b0_mul_componentxUMxa10_and_b1,
         input_times_b0_mul_componentxUMxa9_and_b2,
         input_times_b0_mul_componentxUMxsum_layer1_127732368_127722048_127723952,
         input_times_b0_mul_componentxUMxa8_and_b3,
         input_times_b0_mul_componentxUMxa7_and_b4,
         input_times_b0_mul_componentxUMxa6_and_b5,
         input_times_b0_mul_componentxUMxsum_layer1_127673344_127675248_127730464,
         input_times_b0_mul_componentxUMxa5_and_b6,
         input_times_b0_mul_componentxUMxa4_and_b7,
         input_times_b0_mul_componentxUMxa3_and_b8,
         input_times_b0_mul_componentxUMxsum_layer1_127831344_127845600_127847504,
         input_times_b0_mul_componentxUMxa2_and_b9,
         input_times_b0_mul_componentxUMxa1_and_b10,
         input_times_b0_mul_componentxUMxa0_and_b11,
         input_times_b0_mul_componentxUMxcarry_layer1_127635696_127637600,
         input_times_b0_mul_componentxUMxsum_layer1_127635696_127637600,
         input_times_b0_mul_componentxUMxa10_and_b0,
         input_times_b0_mul_componentxUMxa9_and_b1,
         input_times_b0_mul_componentxUMxsum_layer1_127732256_127721936_127723840,
         input_times_b0_mul_componentxUMxa8_and_b2,
         input_times_b0_mul_componentxUMxa7_and_b3,
         input_times_b0_mul_componentxUMxa6_and_b4,
         input_times_b0_mul_componentxUMxsum_layer1_127673232_127675136_127730352,
         input_times_b0_mul_componentxUMxa5_and_b5,
         input_times_b0_mul_componentxUMxa4_and_b6,
         input_times_b0_mul_componentxUMxa3_and_b7,
         input_times_b0_mul_componentxUMxsum_layer1_127831232_127845488_127847392,
         input_times_b0_mul_componentxUMxa2_and_b8,
         input_times_b0_mul_componentxUMxa1_and_b9,
         input_times_b0_mul_componentxUMxa0_and_b10,
         input_times_b0_mul_componentxUMxsum_layer1_127732144_127721824_127723728,
         input_times_b0_mul_componentxUMxa8_and_b1,
         input_times_b0_mul_componentxUMxa7_and_b2,
         input_times_b0_mul_componentxUMxa6_and_b3,
         input_times_b0_mul_componentxUMxsum_layer1_127673120_127675024_127730240,
         input_times_b0_mul_componentxUMxa5_and_b4,
         input_times_b0_mul_componentxUMxa4_and_b5,
         input_times_b0_mul_componentxUMxa3_and_b6,
         input_times_b0_mul_componentxUMxsum_layer1_127831120_127845376_127847280,
         input_times_b0_mul_componentxUMxa2_and_b7,
         input_times_b0_mul_componentxUMxa1_and_b8,
         input_times_b0_mul_componentxUMxa0_and_b9,
         input_times_b0_mul_componentxUMxsum_layer1_127732032_127721712_127723616,
         input_times_b0_mul_componentxUMxa8_and_b0,
         input_times_b0_mul_componentxUMxa7_and_b1,
         input_times_b0_mul_componentxUMxa6_and_b2,
         input_times_b0_mul_componentxUMxsum_layer1_127673008_127674912_127730128,
         input_times_b0_mul_componentxUMxa5_and_b3,
         input_times_b0_mul_componentxUMxa4_and_b4,
         input_times_b0_mul_componentxUMxa3_and_b5,
         input_times_b0_mul_componentxUMxsum_layer1_127831008_127845264_127847168,
         input_times_b0_mul_componentxUMxa2_and_b6,
         input_times_b0_mul_componentxUMxa1_and_b7,
         input_times_b0_mul_componentxUMxa0_and_b8,
         input_times_b0_mul_componentxUMxcarry_layer1_127731920_127721600,
         input_times_b0_mul_componentxUMxsum_layer1_127731920_127721600,
         input_times_b0_mul_componentxUMxa7_and_b0,
         input_times_b0_mul_componentxUMxa6_and_b1,
         input_times_b0_mul_componentxUMxsum_layer1_127672896_127674800_127730016,
         input_times_b0_mul_componentxUMxa5_and_b2,
         input_times_b0_mul_componentxUMxa4_and_b3,
         input_times_b0_mul_componentxUMxa3_and_b4,
         input_times_b0_mul_componentxUMxsum_layer1_127830896_127845152_127847056,
         input_times_b0_mul_componentxUMxa2_and_b5,
         input_times_b0_mul_componentxUMxa1_and_b6,
         input_times_b0_mul_componentxUMxa0_and_b7,
         input_times_b0_mul_componentxUMxsum_layer1_127672784_127674688_127729904,
         input_times_b0_mul_componentxUMxa5_and_b1,
         input_times_b0_mul_componentxUMxa4_and_b2,
         input_times_b0_mul_componentxUMxa3_and_b3,
         input_times_b0_mul_componentxUMxsum_layer1_127830784_127845040_127846944,
         input_times_b0_mul_componentxUMxa2_and_b4,
         input_times_b0_mul_componentxUMxa1_and_b5,
         input_times_b0_mul_componentxUMxa0_and_b6,
         input_times_b0_mul_componentxUMxsum_layer1_127672672_127674576_127729792,
         input_times_b0_mul_componentxUMxa5_and_b0,
         input_times_b0_mul_componentxUMxa4_and_b1,
         input_times_b0_mul_componentxUMxa3_and_b2,
         input_times_b0_mul_componentxUMxsum_layer1_127830672_127844928_127846832,
         input_times_b0_mul_componentxUMxa2_and_b3,
         input_times_b0_mul_componentxUMxa1_and_b4,
         input_times_b0_mul_componentxUMxa0_and_b5,
         input_times_b0_mul_componentxUMxcarry_layer1_127672560_127674464,
         input_times_b0_mul_componentxUMxsum_layer1_127672560_127674464,
         input_times_b0_mul_componentxUMxa4_and_b0,
         input_times_b0_mul_componentxUMxa3_and_b1,
         input_times_b0_mul_componentxUMxsum_layer1_127830560_127844816_127846720,
         input_times_b0_mul_componentxUMxa2_and_b2,
         input_times_b0_mul_componentxUMxa1_and_b3,
         input_times_b0_mul_componentxUMxa0_and_b4,
         input_times_b0_mul_componentxUMxsum_layer1_127830448_127844704_127846608,
         input_times_b0_mul_componentxUMxa2_and_b1,
         input_times_b0_mul_componentxUMxa1_and_b2,
         input_times_b0_mul_componentxUMxa0_and_b3,
         input_times_b0_mul_componentxUMxsum_layer1_127830336_127844592_127846496,
         input_times_b0_mul_componentxUMxa2_and_b0,
         input_times_b0_mul_componentxUMxa1_and_b1,
         input_times_b0_mul_componentxUMxa0_and_b2,
         input_times_b0_mul_componentxUMxcarry_layer1_127830168_127844480,
         input_times_b0_mul_componentxUMxa1_and_b0,
         input_times_b0_mul_componentxUMxa0_and_b1,
         input_times_b0_div_componentxUDxn19,
         input_times_b0_div_componentxUDxn18,
         input_times_b0_div_componentxUDxn17,
         input_times_b0_div_componentxUDxn16,
         input_times_b0_div_componentxUDxn15,
         input_times_b0_div_componentxUDxn14,
         input_times_b0_div_componentxUDxn13,
         input_times_b0_div_componentxUDxn12,
         input_times_b0_div_componentxUDxn11,
         input_times_b0_div_componentxUDxn10,
         input_times_b0_div_componentxUDxn9,
         input_times_b0_div_componentxUDxn8,
         input_times_b0_div_componentxUDxn7,
         input_times_b0_div_componentxUDxn6,
         input_times_b0_div_componentxUDxn5,
         input_times_b0_div_componentxUDxn4,
         input_times_b0_div_componentxUDxn3,
         input_times_b0_div_componentxUDxn1,
         input_times_b0_div_componentxUDxis_less_than,
         input_times_b0_div_componentxUDxcentral_parallel_output_0,
         input_times_b0_div_componentxUDxcentral_parallel_output_1,
         input_times_b0_div_componentxUDxcentral_parallel_output_2,
         input_times_b0_div_componentxUDxcentral_parallel_output_3,
         input_times_b0_div_componentxUDxcentral_parallel_output_4,
         input_times_b0_div_componentxUDxcentral_parallel_output_5,
         input_times_b0_div_componentxUDxcentral_parallel_output_6,
         input_times_b0_div_componentxUDxcentral_parallel_output_7,
         input_times_b0_div_componentxUDxcentral_parallel_output_8,
         input_times_b0_div_componentxUDxcentral_parallel_output_9,
         input_times_b0_div_componentxUDxcentral_parallel_output_10,
         input_times_b0_div_componentxUDxcentral_parallel_output_11,
         input_times_b0_div_componentxUDxcentral_parallel_output_12,
         input_times_b0_div_componentxUDxcentral_parallel_output_13,
         input_times_b0_div_componentxUDxcentral_parallel_output_14,
         input_times_b0_div_componentxUDxcentral_parallel_output_15,
         input_times_b0_div_componentxUDxcentral_parallel_output_16,
         input_times_b0_div_componentxUDxcentral_parallel_output_17,
         input_times_b0_div_componentxUDxshifted_substraction_result_0,
         input_times_b0_mul_componentxUMxFA_127826296_127826240xn3,
         input_times_b0_mul_componentxUMxFA_127826296_127826240xn2,
         input_times_b0_mul_componentxUMxAdder_finalxn629,
         input_times_b0_mul_componentxUMxAdder_finalxn628,
         input_times_b0_mul_componentxUMxAdder_finalxn607,
         input_times_b0_mul_componentxUMxAdder_finalxn606,
         input_times_b0_mul_componentxUMxAdder_finalxn585,
         input_times_b0_mul_componentxUMxAdder_finalxn584,
         input_times_b0_mul_componentxUMxAdder_finalxn563,
         input_times_b0_mul_componentxUMxAdder_finalxn562,
         input_times_b0_mul_componentxUMxAdder_finalxn541,
         input_times_b0_mul_componentxUMxAdder_finalxn540,
         input_times_b0_mul_componentxUMxAdder_finalxn519,
         input_times_b0_mul_componentxUMxAdder_finalxn518,
         input_times_b0_mul_componentxUMxAdder_finalxn497,
         input_times_b0_mul_componentxUMxAdder_finalxn496,
         input_times_b0_mul_componentxUMxAdder_finalxn475,
         input_times_b0_mul_componentxUMxAdder_finalxn474,
         input_times_b0_mul_componentxUMxAdder_finalxn47,
         input_times_b0_mul_componentxUMxAdder_finalxn25,
         input_times_b0_mul_componentxUMxAdder_finalxn24,
         input_times_b0_mul_componentxUMxAdder_finalxn3,
         input_times_b0_mul_componentxUMxAdder_finalxn2,
         input_times_b0_div_componentxUDxinput_containerxn40,
         input_times_b0_div_componentxUDxinput_containerxn38,
         input_times_b0_div_componentxUDxinput_containerxn37,
         input_times_b0_div_componentxUDxinput_containerxn36,
         input_times_b0_div_componentxUDxinput_containerxn35,
         input_times_b0_div_componentxUDxinput_containerxn34,
         input_times_b0_div_componentxUDxinput_containerxn33,
         input_times_b0_div_componentxUDxinput_containerxn32,
         input_times_b0_div_componentxUDxinput_containerxn31,
         input_times_b0_div_componentxUDxinput_containerxn30,
         input_times_b0_div_componentxUDxinput_containerxn29,
         input_times_b0_div_componentxUDxinput_containerxn28,
         input_times_b0_div_componentxUDxinput_containerxn27,
         input_times_b0_div_componentxUDxinput_containerxn26,
         input_times_b0_div_componentxUDxinput_containerxn25,
         input_times_b0_div_componentxUDxinput_containerxn24,
         input_times_b0_div_componentxUDxinput_containerxn23,
         input_times_b0_div_componentxUDxinput_containerxn22,
         input_times_b0_div_componentxUDxinput_containerxn21,
         input_times_b0_div_componentxUDxinput_containerxn20,
         input_times_b0_div_componentxUDxinput_containerxn19,
         input_times_b0_div_componentxUDxinput_containerxn18,
         input_times_b0_div_componentxUDxinput_containerxn17,
         input_times_b0_div_componentxUDxinput_containerxn16,
         input_times_b0_div_componentxUDxinput_containerxn15,
         input_times_b0_div_componentxUDxinput_containerxn14,
         input_times_b0_div_componentxUDxinput_containerxn13,
         input_times_b0_div_componentxUDxinput_containerxn12,
         input_times_b0_div_componentxUDxinput_containerxn11,
         input_times_b0_div_componentxUDxinput_containerxn10,
         input_times_b0_div_componentxUDxinput_containerxn9,
         input_times_b0_div_componentxUDxinput_containerxn8,
         input_times_b0_div_componentxUDxinput_containerxn7,
         input_times_b0_div_componentxUDxinput_containerxn6,
         input_times_b0_div_componentxUDxinput_containerxn5,
         input_times_b0_div_componentxUDxinput_containerxn3,
         input_times_b0_div_componentxUDxinput_containerxn2,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_0,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_1,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_2,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_3,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_4,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_5,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_6,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_7,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_8,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_9,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_10,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_11,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_12,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_13,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_14,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_15,
         input_times_b0_div_componentxUDxinput_containerxparallel_out_16,
         input_times_b0_div_componentxUDxinverter_for_substractionxn18,
         input_times_b0_div_componentxUDxinverter_for_substractionxn16,
         input_times_b0_div_componentxUDxinverter_for_substractionxn14,
         input_times_b0_div_componentxUDxinverter_for_substractionxn12,
         input_times_b0_div_componentxUDxinverter_for_substractionxn9,
         input_times_b0_div_componentxUDxinverter_for_substractionxn8,
         input_times_b0_div_componentxUDxinverter_for_substractionxn6,
         input_times_b0_div_componentxUDxinverter_for_substractionxn4,
         input_times_b0_div_componentxUDxinverter_for_substractionxn2,
         input_times_b0_div_componentxUDxactually_substractsxn36,
         input_times_b0_div_componentxUDxactually_substractsxn35,
         input_times_b0_div_componentxUDxactually_substractsxn34,
         input_times_b0_div_componentxUDxactually_substractsxn33,
         input_times_b0_div_componentxUDxactually_substractsxn32,
         input_times_b0_div_componentxUDxactually_substractsxn31,
         input_times_b0_div_componentxUDxactually_substractsxn30,
         input_times_b0_div_componentxUDxactually_substractsxn29,
         input_times_b0_div_componentxUDxactually_substractsxn28,
         input_times_b0_div_componentxUDxactually_substractsxn27,
         input_times_b0_div_componentxUDxactually_substractsxn26,
         input_times_b0_div_componentxUDxactually_substractsxn25,
         input_times_b0_div_componentxUDxactually_substractsxn24,
         input_times_b0_div_componentxUDxactually_substractsxn23,
         input_times_b0_div_componentxUDxactually_substractsxn18,
         input_times_b0_div_componentxUDxactually_substractsxn17,
         input_times_b0_div_componentxUDxactually_substractsxn16,
         input_times_b0_div_componentxUDxactually_substractsxn15,
         input_times_b0_div_componentxUDxactually_substractsxn14,
         input_times_b0_div_componentxUDxactually_substractsxn13,
         input_times_b0_div_componentxUDxactually_substractsxn12,
         input_times_b0_div_componentxUDxactually_substractsxn11,
         input_times_b0_div_componentxUDxactually_substractsxn10,
         input_times_b0_div_componentxUDxactually_substractsxn9,
         input_times_b0_div_componentxUDxactually_substractsxn8,
         input_times_b0_div_componentxUDxactually_substractsxn7,
         input_times_b0_div_componentxUDxactually_substractsxn6,
         input_times_b0_div_componentxUDxactually_substractsxn5,
         input_times_b0_div_componentxUDxactually_substractsxn4,
         input_times_b0_div_componentxUDxactually_substractsxn3,
         input_times_b0_div_componentxUDxactually_substractsxn2,
         input_times_b0_div_componentxUDxactually_substractsxn1,
         output_p2_times_a2_mul_componentxunsigned_output_8,
         output_p2_times_a2_mul_componentxunsigned_output_9,
         output_p2_times_a2_mul_componentxunsigned_output_10,
         output_p2_times_a2_mul_componentxunsigned_output_11,
         output_p2_times_a2_mul_componentxunsigned_output_12,
         output_p2_times_a2_mul_componentxunsigned_output_13,
         output_p2_times_a2_mul_componentxunsigned_output_14,
         output_p2_times_a2_mul_componentxunsigned_output_15,
         output_p2_times_a2_mul_componentxunsigned_output_16,
         output_p2_times_a2_mul_componentxunsigned_output_17,
         output_p2_times_a2_mul_componentxinput_B_inverted_1_,
         output_p2_times_a2_mul_componentxinput_B_inverted_2_,
         output_p2_times_a2_mul_componentxinput_B_inverted_3_,
         output_p2_times_a2_mul_componentxinput_B_inverted_4_,
         output_p2_times_a2_mul_componentxinput_B_inverted_5_,
         output_p2_times_a2_mul_componentxinput_B_inverted_6_,
         output_p2_times_a2_mul_componentxinput_B_inverted_7_,
         output_p2_times_a2_mul_componentxinput_B_inverted_8_,
         output_p2_times_a2_mul_componentxinput_B_inverted_9_,
         output_p2_times_a2_mul_componentxinput_B_inverted_10_,
         output_p2_times_a2_mul_componentxinput_B_inverted_11_,
         output_p2_times_a2_mul_componentxinput_B_inverted_12_,
         output_p2_times_a2_mul_componentxinput_B_inverted_13_,
         output_p2_times_a2_mul_componentxinput_B_inverted_14_,
         output_p2_times_a2_mul_componentxinput_B_inverted_15_,
         output_p2_times_a2_mul_componentxinput_B_inverted_16_,
         output_p2_times_a2_mul_componentxinput_B_inverted_17_,
         output_p1_times_a1_mul_componentxunsigned_output_8,
         output_p1_times_a1_mul_componentxunsigned_output_9,
         output_p1_times_a1_mul_componentxunsigned_output_10,
         output_p1_times_a1_mul_componentxunsigned_output_11,
         output_p1_times_a1_mul_componentxunsigned_output_12,
         output_p1_times_a1_mul_componentxunsigned_output_13,
         output_p1_times_a1_mul_componentxunsigned_output_14,
         output_p1_times_a1_mul_componentxunsigned_output_15,
         output_p1_times_a1_mul_componentxunsigned_output_16,
         output_p1_times_a1_mul_componentxunsigned_output_17,
         output_p1_times_a1_mul_componentxinput_B_inverted_1_,
         output_p1_times_a1_mul_componentxinput_B_inverted_2_,
         output_p1_times_a1_mul_componentxinput_B_inverted_3_,
         output_p1_times_a1_mul_componentxinput_B_inverted_4_,
         output_p1_times_a1_mul_componentxinput_B_inverted_5_,
         output_p1_times_a1_mul_componentxinput_B_inverted_6_,
         output_p1_times_a1_mul_componentxinput_B_inverted_7_,
         output_p1_times_a1_mul_componentxinput_B_inverted_8_,
         output_p1_times_a1_mul_componentxinput_B_inverted_9_,
         output_p1_times_a1_mul_componentxinput_B_inverted_10_,
         output_p1_times_a1_mul_componentxinput_B_inverted_11_,
         output_p1_times_a1_mul_componentxinput_B_inverted_12_,
         output_p1_times_a1_mul_componentxinput_B_inverted_13_,
         output_p1_times_a1_mul_componentxinput_B_inverted_14_,
         output_p1_times_a1_mul_componentxinput_B_inverted_15_,
         output_p1_times_a1_mul_componentxinput_B_inverted_16_,
         output_p1_times_a1_mul_componentxinput_B_inverted_17_,
         output_p1_times_a1_mul_componentxinput_A_inverted_1_,
         output_p1_times_a1_mul_componentxinput_A_inverted_2_,
         output_p1_times_a1_mul_componentxinput_A_inverted_3_,
         output_p1_times_a1_mul_componentxinput_A_inverted_4_,
         output_p1_times_a1_mul_componentxinput_A_inverted_5_,
         output_p1_times_a1_mul_componentxinput_A_inverted_6_,
         output_p1_times_a1_mul_componentxinput_A_inverted_7_,
         output_p1_times_a1_mul_componentxinput_A_inverted_8_,
         output_p1_times_a1_mul_componentxinput_A_inverted_9_,
         output_p1_times_a1_mul_componentxinput_A_inverted_10_,
         output_p1_times_a1_mul_componentxinput_A_inverted_11_,
         output_p1_times_a1_mul_componentxinput_A_inverted_12_,
         output_p1_times_a1_mul_componentxinput_A_inverted_13_,
         output_p1_times_a1_mul_componentxinput_A_inverted_14_,
         output_p1_times_a1_mul_componentxinput_A_inverted_15_,
         output_p1_times_a1_mul_componentxinput_A_inverted_16_,
         output_p1_times_a1_mul_componentxinput_A_inverted_17_,
         input_p2_times_b2_mul_componentxunsigned_output_8,
         input_p2_times_b2_mul_componentxunsigned_output_9,
         input_p2_times_b2_mul_componentxunsigned_output_10,
         input_p2_times_b2_mul_componentxunsigned_output_11,
         input_p2_times_b2_mul_componentxunsigned_output_12,
         input_p2_times_b2_mul_componentxunsigned_output_13,
         input_p2_times_b2_mul_componentxunsigned_output_14,
         input_p2_times_b2_mul_componentxunsigned_output_15,
         input_p2_times_b2_mul_componentxunsigned_output_16,
         input_p2_times_b2_mul_componentxunsigned_output_17,
         input_p2_times_b2_mul_componentxinput_B_inverted_1_,
         input_p2_times_b2_mul_componentxinput_B_inverted_2_,
         input_p2_times_b2_mul_componentxinput_B_inverted_3_,
         input_p2_times_b2_mul_componentxinput_B_inverted_4_,
         input_p2_times_b2_mul_componentxinput_B_inverted_5_,
         input_p2_times_b2_mul_componentxinput_B_inverted_6_,
         input_p2_times_b2_mul_componentxinput_B_inverted_7_,
         input_p2_times_b2_mul_componentxinput_B_inverted_8_,
         input_p2_times_b2_mul_componentxinput_B_inverted_9_,
         input_p2_times_b2_mul_componentxinput_B_inverted_10_,
         input_p2_times_b2_mul_componentxinput_B_inverted_11_,
         input_p2_times_b2_mul_componentxinput_B_inverted_12_,
         input_p2_times_b2_mul_componentxinput_B_inverted_13_,
         input_p2_times_b2_mul_componentxinput_B_inverted_14_,
         input_p2_times_b2_mul_componentxinput_B_inverted_15_,
         input_p2_times_b2_mul_componentxinput_B_inverted_16_,
         input_p2_times_b2_mul_componentxinput_B_inverted_17_,
         input_p1_times_b1_mul_componentxunsigned_output_8,
         input_p1_times_b1_mul_componentxunsigned_output_9,
         input_p1_times_b1_mul_componentxunsigned_output_10,
         input_p1_times_b1_mul_componentxunsigned_output_11,
         input_p1_times_b1_mul_componentxunsigned_output_12,
         input_p1_times_b1_mul_componentxunsigned_output_13,
         input_p1_times_b1_mul_componentxunsigned_output_14,
         input_p1_times_b1_mul_componentxunsigned_output_15,
         input_p1_times_b1_mul_componentxunsigned_output_16,
         input_p1_times_b1_mul_componentxunsigned_output_17,
         input_p1_times_b1_mul_componentxinput_B_inverted_1_,
         input_p1_times_b1_mul_componentxinput_B_inverted_2_,
         input_p1_times_b1_mul_componentxinput_B_inverted_3_,
         input_p1_times_b1_mul_componentxinput_B_inverted_4_,
         input_p1_times_b1_mul_componentxinput_B_inverted_5_,
         input_p1_times_b1_mul_componentxinput_B_inverted_6_,
         input_p1_times_b1_mul_componentxinput_B_inverted_7_,
         input_p1_times_b1_mul_componentxinput_B_inverted_8_,
         input_p1_times_b1_mul_componentxinput_B_inverted_9_,
         input_p1_times_b1_mul_componentxinput_B_inverted_10_,
         input_p1_times_b1_mul_componentxinput_B_inverted_11_,
         input_p1_times_b1_mul_componentxinput_B_inverted_12_,
         input_p1_times_b1_mul_componentxinput_B_inverted_13_,
         input_p1_times_b1_mul_componentxinput_B_inverted_14_,
         input_p1_times_b1_mul_componentxinput_B_inverted_15_,
         input_p1_times_b1_mul_componentxinput_B_inverted_16_,
         input_p1_times_b1_mul_componentxinput_B_inverted_17_,
         output_p2_times_a2_div_componentxoutput_sign_gated,
         output_p2_times_a2_div_componentxoutput_sign_gated_prev,
         output_p2_times_a2_div_componentxunsigned_B_17,
         output_p2_times_a2_div_componentxunsigned_A_17,
         output_p2_times_a2_div_componentxunsigned_output_1,
         output_p2_times_a2_div_componentxunsigned_output_2,
         output_p2_times_a2_div_componentxunsigned_output_3,
         output_p2_times_a2_div_componentxunsigned_output_4,
         output_p2_times_a2_div_componentxunsigned_output_5,
         output_p2_times_a2_div_componentxunsigned_output_6,
         output_p2_times_a2_div_componentxunsigned_output_7,
         output_p2_times_a2_div_componentxunsigned_output_8,
         output_p2_times_a2_div_componentxunsigned_output_9,
         output_p2_times_a2_div_componentxunsigned_output_10,
         output_p2_times_a2_div_componentxunsigned_output_11,
         output_p2_times_a2_div_componentxunsigned_output_12,
         output_p2_times_a2_div_componentxunsigned_output_13,
         output_p2_times_a2_div_componentxunsigned_output_14,
         output_p2_times_a2_div_componentxunsigned_output_15,
         output_p2_times_a2_div_componentxunsigned_output_16,
         output_p2_times_a2_div_componentxunsigned_output_17,
         output_p2_times_a2_div_componentxinput_B_inverted_1_,
         output_p2_times_a2_div_componentxinput_B_inverted_2_,
         output_p2_times_a2_div_componentxinput_B_inverted_3_,
         output_p2_times_a2_div_componentxinput_B_inverted_4_,
         output_p2_times_a2_div_componentxinput_B_inverted_5_,
         output_p2_times_a2_div_componentxinput_B_inverted_6_,
         output_p2_times_a2_div_componentxinput_B_inverted_7_,
         output_p2_times_a2_div_componentxinput_B_inverted_8_,
         output_p2_times_a2_div_componentxinput_B_inverted_9_,
         output_p2_times_a2_div_componentxinput_B_inverted_10_,
         output_p2_times_a2_div_componentxinput_B_inverted_11_,
         output_p2_times_a2_div_componentxinput_B_inverted_12_,
         output_p2_times_a2_div_componentxinput_B_inverted_13_,
         output_p2_times_a2_div_componentxinput_B_inverted_14_,
         output_p2_times_a2_div_componentxinput_B_inverted_15_,
         output_p2_times_a2_div_componentxinput_B_inverted_16_,
         output_p2_times_a2_div_componentxinput_B_inverted_17_,
         output_p1_times_a1_div_componentxoutput_sign_gated,
         output_p1_times_a1_div_componentxoutput_ready_signal,
         output_p1_times_a1_div_componentxunsigned_B_17,
         output_p1_times_a1_div_componentxunsigned_A_17,
         output_p1_times_a1_div_componentxunsigned_output_1,
         output_p1_times_a1_div_componentxunsigned_output_2,
         output_p1_times_a1_div_componentxunsigned_output_3,
         output_p1_times_a1_div_componentxunsigned_output_4,
         output_p1_times_a1_div_componentxunsigned_output_5,
         output_p1_times_a1_div_componentxunsigned_output_6,
         output_p1_times_a1_div_componentxunsigned_output_7,
         output_p1_times_a1_div_componentxunsigned_output_8,
         output_p1_times_a1_div_componentxunsigned_output_9,
         output_p1_times_a1_div_componentxunsigned_output_10,
         output_p1_times_a1_div_componentxunsigned_output_11,
         output_p1_times_a1_div_componentxunsigned_output_12,
         output_p1_times_a1_div_componentxunsigned_output_13,
         output_p1_times_a1_div_componentxunsigned_output_14,
         output_p1_times_a1_div_componentxunsigned_output_15,
         output_p1_times_a1_div_componentxunsigned_output_16,
         output_p1_times_a1_div_componentxunsigned_output_17,
         output_p1_times_a1_div_componentxinput_B_inverted_1_,
         output_p1_times_a1_div_componentxinput_B_inverted_2_,
         output_p1_times_a1_div_componentxinput_B_inverted_3_,
         output_p1_times_a1_div_componentxinput_B_inverted_4_,
         output_p1_times_a1_div_componentxinput_B_inverted_5_,
         output_p1_times_a1_div_componentxinput_B_inverted_6_,
         output_p1_times_a1_div_componentxinput_B_inverted_7_,
         output_p1_times_a1_div_componentxinput_B_inverted_8_,
         output_p1_times_a1_div_componentxinput_B_inverted_9_,
         output_p1_times_a1_div_componentxinput_B_inverted_10_,
         output_p1_times_a1_div_componentxinput_B_inverted_11_,
         output_p1_times_a1_div_componentxinput_B_inverted_12_,
         output_p1_times_a1_div_componentxinput_B_inverted_13_,
         output_p1_times_a1_div_componentxinput_B_inverted_14_,
         output_p1_times_a1_div_componentxinput_B_inverted_15_,
         output_p1_times_a1_div_componentxinput_B_inverted_16_,
         output_p1_times_a1_div_componentxinput_B_inverted_17_,
         input_p2_times_b2_div_componentxoutput_sign_gated,
         input_p2_times_b2_div_componentxoutput_sign_gated_prev,
         input_p2_times_b2_div_componentxoutput_ready_signal,
         input_p2_times_b2_div_componentxunsigned_B_17,
         input_p2_times_b2_div_componentxunsigned_A_17,
         input_p2_times_b2_div_componentxunsigned_output_1,
         input_p2_times_b2_div_componentxunsigned_output_2,
         input_p2_times_b2_div_componentxunsigned_output_3,
         input_p2_times_b2_div_componentxunsigned_output_4,
         input_p2_times_b2_div_componentxunsigned_output_5,
         input_p2_times_b2_div_componentxunsigned_output_6,
         input_p2_times_b2_div_componentxunsigned_output_7,
         input_p2_times_b2_div_componentxunsigned_output_8,
         input_p2_times_b2_div_componentxunsigned_output_9,
         input_p2_times_b2_div_componentxunsigned_output_10,
         input_p2_times_b2_div_componentxunsigned_output_11,
         input_p2_times_b2_div_componentxunsigned_output_12,
         input_p2_times_b2_div_componentxunsigned_output_13,
         input_p2_times_b2_div_componentxunsigned_output_14,
         input_p2_times_b2_div_componentxunsigned_output_15,
         input_p2_times_b2_div_componentxunsigned_output_16,
         input_p2_times_b2_div_componentxunsigned_output_17,
         input_p2_times_b2_div_componentxinput_B_inverted_1_,
         input_p2_times_b2_div_componentxinput_B_inverted_2_,
         input_p2_times_b2_div_componentxinput_B_inverted_3_,
         input_p2_times_b2_div_componentxinput_B_inverted_4_,
         input_p2_times_b2_div_componentxinput_B_inverted_5_,
         input_p2_times_b2_div_componentxinput_B_inverted_6_,
         input_p2_times_b2_div_componentxinput_B_inverted_7_,
         input_p2_times_b2_div_componentxinput_B_inverted_8_,
         input_p2_times_b2_div_componentxinput_B_inverted_9_,
         input_p2_times_b2_div_componentxinput_B_inverted_10_,
         input_p2_times_b2_div_componentxinput_B_inverted_11_,
         input_p2_times_b2_div_componentxinput_B_inverted_12_,
         input_p2_times_b2_div_componentxinput_B_inverted_13_,
         input_p2_times_b2_div_componentxinput_B_inverted_14_,
         input_p2_times_b2_div_componentxinput_B_inverted_15_,
         input_p2_times_b2_div_componentxinput_B_inverted_16_,
         input_p2_times_b2_div_componentxinput_B_inverted_17_,
         input_p1_times_b1_div_componentxoutput_sign_gated,
         input_p1_times_b1_div_componentxoutput_sign_gated_prev,
         input_p1_times_b1_div_componentxoutput_ready_signal,
         input_p1_times_b1_div_componentxunsigned_B_17,
         input_p1_times_b1_div_componentxunsigned_A_17,
         input_p1_times_b1_div_componentxunsigned_output_1,
         input_p1_times_b1_div_componentxunsigned_output_2,
         input_p1_times_b1_div_componentxunsigned_output_3,
         input_p1_times_b1_div_componentxunsigned_output_4,
         input_p1_times_b1_div_componentxunsigned_output_5,
         input_p1_times_b1_div_componentxunsigned_output_6,
         input_p1_times_b1_div_componentxunsigned_output_7,
         input_p1_times_b1_div_componentxunsigned_output_8,
         input_p1_times_b1_div_componentxunsigned_output_9,
         input_p1_times_b1_div_componentxunsigned_output_10,
         input_p1_times_b1_div_componentxunsigned_output_11,
         input_p1_times_b1_div_componentxunsigned_output_12,
         input_p1_times_b1_div_componentxunsigned_output_13,
         input_p1_times_b1_div_componentxunsigned_output_14,
         input_p1_times_b1_div_componentxunsigned_output_15,
         input_p1_times_b1_div_componentxunsigned_output_16,
         input_p1_times_b1_div_componentxunsigned_output_17,
         input_p1_times_b1_div_componentxinput_B_inverted_1_,
         input_p1_times_b1_div_componentxinput_B_inverted_2_,
         input_p1_times_b1_div_componentxinput_B_inverted_3_,
         input_p1_times_b1_div_componentxinput_B_inverted_4_,
         input_p1_times_b1_div_componentxinput_B_inverted_5_,
         input_p1_times_b1_div_componentxinput_B_inverted_6_,
         input_p1_times_b1_div_componentxinput_B_inverted_7_,
         input_p1_times_b1_div_componentxinput_B_inverted_8_,
         input_p1_times_b1_div_componentxinput_B_inverted_9_,
         input_p1_times_b1_div_componentxinput_B_inverted_10_,
         input_p1_times_b1_div_componentxinput_B_inverted_11_,
         input_p1_times_b1_div_componentxinput_B_inverted_12_,
         input_p1_times_b1_div_componentxinput_B_inverted_13_,
         input_p1_times_b1_div_componentxinput_B_inverted_14_,
         input_p1_times_b1_div_componentxinput_B_inverted_15_,
         input_p1_times_b1_div_componentxinput_B_inverted_16_,
         input_p1_times_b1_div_componentxinput_B_inverted_17_,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128315744_128315968_128316136,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128315464_128315632_128315800,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128220800_128221024_128221136,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128220688_128220856_128220968,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128126256_128220520_128220744,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128125920_128220352_128220576,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128125584_128220184_128220408,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128125248_128219960_128220240,
         output_p2_times_a2_mul_componentxUMxcarry_layer5_128219792_128220016,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128219792_128220016,
         output_p2_times_a2_mul_componentxUMxcarry_layer5_128219624_128219848,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128219624_128219848,
         output_p2_times_a2_mul_componentxUMxcarry_layer5_128219456_128219680,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128219456_128219680,
         output_p2_times_a2_mul_componentxUMxcarry_layer5_128219288_128219512,
         output_p2_times_a2_mul_componentxUMxsum_layer5_128219288_128219512,
         output_p2_times_a2_mul_componentxUMxcarry_layer5_128219120_128219344,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128238312_128238424_128238592,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128237752_128237976_128238144,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128237920_128238088,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128126760_128237640_128237808,
         output_p2_times_a2_mul_componentxUMxcarry_layer4_128126816_128126928,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128126816_128126928,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128263168_128126424_128126648,
         output_p2_times_a2_mul_componentxUMxcarry_layer4_128126480_128126592,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128126480_128126592,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128262496_128126088_128126312,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128125752_128125976_128126144,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128125416_128125640_128125808,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128125080_128125304_128125472,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128124744_128124968_128125136,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128124632_128124800_128124912,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128247456_128124464_128124688,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128247120_128124240_128124520,
         output_p2_times_a2_mul_componentxUMxcarry_layer4_128124072_128124296,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128124072_128124296,
         output_p2_times_a2_mul_componentxUMxcarry_layer4_128123904_128124128,
         output_p2_times_a2_mul_componentxUMxsum_layer4_128123904_128124128,
         output_p2_times_a2_mul_componentxUMxcarry_layer4_128123792_128123960,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128264344_128264512,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128263896_128264064_128264176,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128263336_128263560_128263728,
         output_p2_times_a2_mul_componentxUMxcarry_layer3_128263672_128263840,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128263672_128263840,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128263224_128263392_128263504,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128262664_128262888_128263056,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128262720_128262832_128263000,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128262216_128262384_128262552,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128249696_128249808_128262328,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128197128_128249304_128249528,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128249360_128249472_128249640,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128248800_128249024_128249192,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128248856_128248968_128249136,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128248296_128248520_128248688,
         output_p2_times_a2_mul_componentxUMxcarry_layer3_128248464_128248632,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128248464_128248632,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128247960_128248184_128248352,
         output_p2_times_a2_mul_componentxUMxcarry_layer3_128248016_128248128,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128248016_128248128,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128222880_128247624_128247848,
         output_p2_times_a2_mul_componentxUMxcarry_layer3_128247680_128247792,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128247680_128247792,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128222208_128247288_128247512,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128246952_128247176_128247344,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128246616_128246840_128247008,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128246504_128246672_128246784,
         output_p2_times_a2_mul_componentxUMxsum_layer3_127827080_128246280_128246560,
         output_p2_times_a2_mul_componentxUMxcarry_layer3_128246112_128246336,
         output_p2_times_a2_mul_componentxUMxsum_layer3_128246112_128246336,
         output_p2_times_a2_mul_componentxUMxcarry_layer3_128246000_128246168,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128199816_128200040_128199984,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128199368_128199480_128199648,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128198864_128199032_128199200,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128198304_128198528_128198696,
         output_p2_times_a2_mul_componentxUMxcarry_layer2_128198976_128199144,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128198976_128199144,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128198472_128198640_128198808,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128198080_128198192_128198360,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128197464_128197688_128197856,
         output_p2_times_a2_mul_componentxUMxcarry_layer2_128198024_128197968,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128198024_128197968,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128197520_128197632_128197800,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128197016_128197240_128197352,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127627392_128196680_128196848,
         output_p2_times_a2_mul_componentxUMxa15_and_b0,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128196792_128196960_128197184,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128224952_128225120_128225232,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128224392_128224616_128224784,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128224728_128224896_128225064,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128224280_128224448_128224560,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128223720_128223944_128224168,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128223888_128224112_128224056,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128223440_128223608_128223776,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127715424_128223048_128223272,
         output_p2_times_a2_mul_componentxUMxa12_and_b0,
         output_p2_times_a2_mul_componentxUMxcarry_layer2_128223384_128223552,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128223384_128223552,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128222936_128223104_128223216,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128222376_128222600_128222768,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128222432_128222544_128222712,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128221872_128222096_128222264,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128221760_128221928_128222040,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127635584_128221368_128221592,
         output_p2_times_a2_mul_componentxUMxa9_and_b0,
         output_p2_times_a2_mul_componentxUMxsum_layer2_128221424_128221536_128221704,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127827584_127827808_128221256,
         output_p2_times_a2_mul_componentxUMxcarry_layer2_127827752_127827920,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127827752_127827920,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127827248_127827472_127827640,
         output_p2_times_a2_mul_componentxUMxcarry_layer2_127827304_127827416,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127827304_127827416,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127731808_127826912_127827136,
         output_p2_times_a2_mul_componentxUMxa6_and_b0,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127826576_127826800_127826968,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127826464_127826632_127826744,
         output_p2_times_a2_mul_componentxUMxsum_layer2_127672448_127826240_127826520,
         output_p2_times_a2_mul_componentxUMxa3_and_b0,
         output_p2_times_a2_mul_componentxUMxcarry_layer2_127826128_127826296,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127627616_127629520_127824000,
         output_p2_times_a2_mul_componentxUMxa17_and_b0,
         output_p2_times_a2_mul_componentxUMxa16_and_b1,
         output_p2_times_a2_mul_componentxUMxa15_and_b2,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127715984_127849024_127850928,
         output_p2_times_a2_mul_componentxUMxa14_and_b3,
         output_p2_times_a2_mul_componentxUMxa13_and_b4,
         output_p2_times_a2_mul_componentxUMxa12_and_b5,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127636480_127638384_127714080,
         output_p2_times_a2_mul_componentxUMxa11_and_b6,
         output_p2_times_a2_mul_componentxUMxa10_and_b7,
         output_p2_times_a2_mul_componentxUMxa9_and_b8,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127733040_127722720_127724624,
         output_p2_times_a2_mul_componentxUMxa8_and_b9,
         output_p2_times_a2_mul_componentxUMxa7_and_b10,
         output_p2_times_a2_mul_componentxUMxa6_and_b11,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127674016_127675920_127731136,
         output_p2_times_a2_mul_componentxUMxa5_and_b12,
         output_p2_times_a2_mul_componentxUMxa4_and_b13,
         output_p2_times_a2_mul_componentxUMxa3_and_b14,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127832016_127846272_127848176,
         output_p2_times_a2_mul_componentxUMxa2_and_b15,
         output_p2_times_a2_mul_componentxUMxa1_and_b16,
         output_p2_times_a2_mul_componentxUMxa0_and_b17,
         output_p2_times_a2_mul_componentxUMxcarry_layer1_127627504_127629408,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127627504_127629408,
         output_p2_times_a2_mul_componentxUMxa16_and_b0,
         output_p2_times_a2_mul_componentxUMxa15_and_b1,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127715872_127848912_127850816,
         output_p2_times_a2_mul_componentxUMxa14_and_b2,
         output_p2_times_a2_mul_componentxUMxa13_and_b3,
         output_p2_times_a2_mul_componentxUMxa12_and_b4,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127636368_127638272_127713968,
         output_p2_times_a2_mul_componentxUMxa11_and_b5,
         output_p2_times_a2_mul_componentxUMxa10_and_b6,
         output_p2_times_a2_mul_componentxUMxa9_and_b7,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732928_127722608_127724512,
         output_p2_times_a2_mul_componentxUMxa8_and_b8,
         output_p2_times_a2_mul_componentxUMxa7_and_b9,
         output_p2_times_a2_mul_componentxUMxa6_and_b10,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673904_127675808_127731024,
         output_p2_times_a2_mul_componentxUMxa5_and_b11,
         output_p2_times_a2_mul_componentxUMxa4_and_b12,
         output_p2_times_a2_mul_componentxUMxa3_and_b13,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831904_127846160_127848064,
         output_p2_times_a2_mul_componentxUMxa2_and_b14,
         output_p2_times_a2_mul_componentxUMxa1_and_b15,
         output_p2_times_a2_mul_componentxUMxa0_and_b16,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127715760_127848800_127850704,
         output_p2_times_a2_mul_componentxUMxa14_and_b1,
         output_p2_times_a2_mul_componentxUMxa13_and_b2,
         output_p2_times_a2_mul_componentxUMxa12_and_b3,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127636256_127638160_127713856,
         output_p2_times_a2_mul_componentxUMxa11_and_b4,
         output_p2_times_a2_mul_componentxUMxa10_and_b5,
         output_p2_times_a2_mul_componentxUMxa9_and_b6,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732816_127722496_127724400,
         output_p2_times_a2_mul_componentxUMxa8_and_b7,
         output_p2_times_a2_mul_componentxUMxa7_and_b8,
         output_p2_times_a2_mul_componentxUMxa6_and_b9,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673792_127675696_127730912,
         output_p2_times_a2_mul_componentxUMxa5_and_b10,
         output_p2_times_a2_mul_componentxUMxa4_and_b11,
         output_p2_times_a2_mul_componentxUMxa3_and_b12,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831792_127846048_127847952,
         output_p2_times_a2_mul_componentxUMxa2_and_b13,
         output_p2_times_a2_mul_componentxUMxa1_and_b14,
         output_p2_times_a2_mul_componentxUMxa0_and_b15,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127715648_127848688_127850592,
         output_p2_times_a2_mul_componentxUMxa14_and_b0,
         output_p2_times_a2_mul_componentxUMxa13_and_b1,
         output_p2_times_a2_mul_componentxUMxa12_and_b2,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127636144_127638048_127713744,
         output_p2_times_a2_mul_componentxUMxa11_and_b3,
         output_p2_times_a2_mul_componentxUMxa10_and_b4,
         output_p2_times_a2_mul_componentxUMxa9_and_b5,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732704_127722384_127724288,
         output_p2_times_a2_mul_componentxUMxa8_and_b6,
         output_p2_times_a2_mul_componentxUMxa7_and_b7,
         output_p2_times_a2_mul_componentxUMxa6_and_b8,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673680_127675584_127730800,
         output_p2_times_a2_mul_componentxUMxa5_and_b9,
         output_p2_times_a2_mul_componentxUMxa4_and_b10,
         output_p2_times_a2_mul_componentxUMxa3_and_b11,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831680_127845936_127847840,
         output_p2_times_a2_mul_componentxUMxa2_and_b12,
         output_p2_times_a2_mul_componentxUMxa1_and_b13,
         output_p2_times_a2_mul_componentxUMxa0_and_b14,
         output_p2_times_a2_mul_componentxUMxcarry_layer1_127715536_127848576,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127715536_127848576,
         output_p2_times_a2_mul_componentxUMxa13_and_b0,
         output_p2_times_a2_mul_componentxUMxa12_and_b1,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127636032_127637936_127713632,
         output_p2_times_a2_mul_componentxUMxa11_and_b2,
         output_p2_times_a2_mul_componentxUMxa10_and_b3,
         output_p2_times_a2_mul_componentxUMxa9_and_b4,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732592_127722272_127724176,
         output_p2_times_a2_mul_componentxUMxa8_and_b5,
         output_p2_times_a2_mul_componentxUMxa7_and_b6,
         output_p2_times_a2_mul_componentxUMxa6_and_b7,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673568_127675472_127730688,
         output_p2_times_a2_mul_componentxUMxa5_and_b8,
         output_p2_times_a2_mul_componentxUMxa4_and_b9,
         output_p2_times_a2_mul_componentxUMxa3_and_b10,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831568_127845824_127847728,
         output_p2_times_a2_mul_componentxUMxa2_and_b11,
         output_p2_times_a2_mul_componentxUMxa1_and_b12,
         output_p2_times_a2_mul_componentxUMxa0_and_b13,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127635920_127637824_127713520,
         output_p2_times_a2_mul_componentxUMxa11_and_b1,
         output_p2_times_a2_mul_componentxUMxa10_and_b2,
         output_p2_times_a2_mul_componentxUMxa9_and_b3,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732480_127722160_127724064,
         output_p2_times_a2_mul_componentxUMxa8_and_b4,
         output_p2_times_a2_mul_componentxUMxa7_and_b5,
         output_p2_times_a2_mul_componentxUMxa6_and_b6,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673456_127675360_127730576,
         output_p2_times_a2_mul_componentxUMxa5_and_b7,
         output_p2_times_a2_mul_componentxUMxa4_and_b8,
         output_p2_times_a2_mul_componentxUMxa3_and_b9,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831456_127845712_127847616,
         output_p2_times_a2_mul_componentxUMxa2_and_b10,
         output_p2_times_a2_mul_componentxUMxa1_and_b11,
         output_p2_times_a2_mul_componentxUMxa0_and_b12,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127635808_127637712_127713408,
         output_p2_times_a2_mul_componentxUMxa11_and_b0,
         output_p2_times_a2_mul_componentxUMxa10_and_b1,
         output_p2_times_a2_mul_componentxUMxa9_and_b2,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732368_127722048_127723952,
         output_p2_times_a2_mul_componentxUMxa8_and_b3,
         output_p2_times_a2_mul_componentxUMxa7_and_b4,
         output_p2_times_a2_mul_componentxUMxa6_and_b5,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673344_127675248_127730464,
         output_p2_times_a2_mul_componentxUMxa5_and_b6,
         output_p2_times_a2_mul_componentxUMxa4_and_b7,
         output_p2_times_a2_mul_componentxUMxa3_and_b8,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831344_127845600_127847504,
         output_p2_times_a2_mul_componentxUMxa2_and_b9,
         output_p2_times_a2_mul_componentxUMxa1_and_b10,
         output_p2_times_a2_mul_componentxUMxa0_and_b11,
         output_p2_times_a2_mul_componentxUMxcarry_layer1_127635696_127637600,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127635696_127637600,
         output_p2_times_a2_mul_componentxUMxa10_and_b0,
         output_p2_times_a2_mul_componentxUMxa9_and_b1,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732256_127721936_127723840,
         output_p2_times_a2_mul_componentxUMxa8_and_b2,
         output_p2_times_a2_mul_componentxUMxa7_and_b3,
         output_p2_times_a2_mul_componentxUMxa6_and_b4,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673232_127675136_127730352,
         output_p2_times_a2_mul_componentxUMxa5_and_b5,
         output_p2_times_a2_mul_componentxUMxa4_and_b6,
         output_p2_times_a2_mul_componentxUMxa3_and_b7,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831232_127845488_127847392,
         output_p2_times_a2_mul_componentxUMxa2_and_b8,
         output_p2_times_a2_mul_componentxUMxa1_and_b9,
         output_p2_times_a2_mul_componentxUMxa0_and_b10,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732144_127721824_127723728,
         output_p2_times_a2_mul_componentxUMxa8_and_b1,
         output_p2_times_a2_mul_componentxUMxa7_and_b2,
         output_p2_times_a2_mul_componentxUMxa6_and_b3,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673120_127675024_127730240,
         output_p2_times_a2_mul_componentxUMxa5_and_b4,
         output_p2_times_a2_mul_componentxUMxa4_and_b5,
         output_p2_times_a2_mul_componentxUMxa3_and_b6,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831120_127845376_127847280,
         output_p2_times_a2_mul_componentxUMxa2_and_b7,
         output_p2_times_a2_mul_componentxUMxa1_and_b8,
         output_p2_times_a2_mul_componentxUMxa0_and_b9,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127732032_127721712_127723616,
         output_p2_times_a2_mul_componentxUMxa8_and_b0,
         output_p2_times_a2_mul_componentxUMxa7_and_b1,
         output_p2_times_a2_mul_componentxUMxa6_and_b2,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127673008_127674912_127730128,
         output_p2_times_a2_mul_componentxUMxa5_and_b3,
         output_p2_times_a2_mul_componentxUMxa4_and_b4,
         output_p2_times_a2_mul_componentxUMxa3_and_b5,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127831008_127845264_127847168,
         output_p2_times_a2_mul_componentxUMxa2_and_b6,
         output_p2_times_a2_mul_componentxUMxa1_and_b7,
         output_p2_times_a2_mul_componentxUMxa0_and_b8,
         output_p2_times_a2_mul_componentxUMxcarry_layer1_127731920_127721600,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127731920_127721600,
         output_p2_times_a2_mul_componentxUMxa7_and_b0,
         output_p2_times_a2_mul_componentxUMxa6_and_b1,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127672896_127674800_127730016,
         output_p2_times_a2_mul_componentxUMxa5_and_b2,
         output_p2_times_a2_mul_componentxUMxa4_and_b3,
         output_p2_times_a2_mul_componentxUMxa3_and_b4,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127830896_127845152_127847056,
         output_p2_times_a2_mul_componentxUMxa2_and_b5,
         output_p2_times_a2_mul_componentxUMxa1_and_b6,
         output_p2_times_a2_mul_componentxUMxa0_and_b7,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127672784_127674688_127729904,
         output_p2_times_a2_mul_componentxUMxa5_and_b1,
         output_p2_times_a2_mul_componentxUMxa4_and_b2,
         output_p2_times_a2_mul_componentxUMxa3_and_b3,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127830784_127845040_127846944,
         output_p2_times_a2_mul_componentxUMxa2_and_b4,
         output_p2_times_a2_mul_componentxUMxa1_and_b5,
         output_p2_times_a2_mul_componentxUMxa0_and_b6,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127672672_127674576_127729792,
         output_p2_times_a2_mul_componentxUMxa5_and_b0,
         output_p2_times_a2_mul_componentxUMxa4_and_b1,
         output_p2_times_a2_mul_componentxUMxa3_and_b2,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127830672_127844928_127846832,
         output_p2_times_a2_mul_componentxUMxa2_and_b3,
         output_p2_times_a2_mul_componentxUMxa1_and_b4,
         output_p2_times_a2_mul_componentxUMxa0_and_b5,
         output_p2_times_a2_mul_componentxUMxcarry_layer1_127672560_127674464,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127672560_127674464,
         output_p2_times_a2_mul_componentxUMxa4_and_b0,
         output_p2_times_a2_mul_componentxUMxa3_and_b1,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127830560_127844816_127846720,
         output_p2_times_a2_mul_componentxUMxa2_and_b2,
         output_p2_times_a2_mul_componentxUMxa1_and_b3,
         output_p2_times_a2_mul_componentxUMxa0_and_b4,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127830448_127844704_127846608,
         output_p2_times_a2_mul_componentxUMxa2_and_b1,
         output_p2_times_a2_mul_componentxUMxa1_and_b2,
         output_p2_times_a2_mul_componentxUMxa0_and_b3,
         output_p2_times_a2_mul_componentxUMxsum_layer1_127830336_127844592_127846496,
         output_p2_times_a2_mul_componentxUMxa2_and_b0,
         output_p2_times_a2_mul_componentxUMxa1_and_b1,
         output_p2_times_a2_mul_componentxUMxa0_and_b2,
         output_p2_times_a2_mul_componentxUMxcarry_layer1_127830168_127844480,
         output_p2_times_a2_mul_componentxUMxa1_and_b0,
         output_p2_times_a2_mul_componentxUMxa0_and_b1,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128315744_128315968_128316136,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128315464_128315632_128315800,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128220800_128221024_128221136,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128220688_128220856_128220968,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128126256_128220520_128220744,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128125920_128220352_128220576,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128125584_128220184_128220408,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128125248_128219960_128220240,
         output_p1_times_a1_mul_componentxUMxcarry_layer5_128219792_128220016,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128219792_128220016,
         output_p1_times_a1_mul_componentxUMxcarry_layer5_128219624_128219848,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128219624_128219848,
         output_p1_times_a1_mul_componentxUMxcarry_layer5_128219456_128219680,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128219456_128219680,
         output_p1_times_a1_mul_componentxUMxcarry_layer5_128219288_128219512,
         output_p1_times_a1_mul_componentxUMxsum_layer5_128219288_128219512,
         output_p1_times_a1_mul_componentxUMxcarry_layer5_128219120_128219344,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128238312_128238424_128238592,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128237752_128237976_128238144,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128237920_128238088,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128126760_128237640_128237808,
         output_p1_times_a1_mul_componentxUMxcarry_layer4_128126816_128126928,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128126816_128126928,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128263168_128126424_128126648,
         output_p1_times_a1_mul_componentxUMxcarry_layer4_128126480_128126592,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128126480_128126592,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128262496_128126088_128126312,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128125752_128125976_128126144,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128125416_128125640_128125808,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128125080_128125304_128125472,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128124744_128124968_128125136,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128124632_128124800_128124912,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128247456_128124464_128124688,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128247120_128124240_128124520,
         output_p1_times_a1_mul_componentxUMxcarry_layer4_128124072_128124296,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128124072_128124296,
         output_p1_times_a1_mul_componentxUMxcarry_layer4_128123904_128124128,
         output_p1_times_a1_mul_componentxUMxsum_layer4_128123904_128124128,
         output_p1_times_a1_mul_componentxUMxcarry_layer4_128123792_128123960,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128264344_128264512,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128263896_128264064_128264176,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128263336_128263560_128263728,
         output_p1_times_a1_mul_componentxUMxcarry_layer3_128263672_128263840,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128263672_128263840,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128263224_128263392_128263504,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128262664_128262888_128263056,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128262720_128262832_128263000,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128262216_128262384_128262552,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128249696_128249808_128262328,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128197128_128249304_128249528,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128249360_128249472_128249640,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128248800_128249024_128249192,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128248856_128248968_128249136,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128248296_128248520_128248688,
         output_p1_times_a1_mul_componentxUMxcarry_layer3_128248464_128248632,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128248464_128248632,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128247960_128248184_128248352,
         output_p1_times_a1_mul_componentxUMxcarry_layer3_128248016_128248128,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128248016_128248128,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128222880_128247624_128247848,
         output_p1_times_a1_mul_componentxUMxcarry_layer3_128247680_128247792,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128247680_128247792,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128222208_128247288_128247512,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128246952_128247176_128247344,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128246616_128246840_128247008,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128246504_128246672_128246784,
         output_p1_times_a1_mul_componentxUMxsum_layer3_127827080_128246280_128246560,
         output_p1_times_a1_mul_componentxUMxcarry_layer3_128246112_128246336,
         output_p1_times_a1_mul_componentxUMxsum_layer3_128246112_128246336,
         output_p1_times_a1_mul_componentxUMxcarry_layer3_128246000_128246168,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128199816_128200040_128199984,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128199368_128199480_128199648,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128198864_128199032_128199200,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128198304_128198528_128198696,
         output_p1_times_a1_mul_componentxUMxcarry_layer2_128198976_128199144,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128198976_128199144,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128198472_128198640_128198808,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128198080_128198192_128198360,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128197464_128197688_128197856,
         output_p1_times_a1_mul_componentxUMxcarry_layer2_128198024_128197968,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128198024_128197968,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128197520_128197632_128197800,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128197016_128197240_128197352,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127627392_128196680_128196848,
         output_p1_times_a1_mul_componentxUMxa15_and_b0,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128196792_128196960_128197184,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128224952_128225120_128225232,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128224392_128224616_128224784,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128224728_128224896_128225064,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128224280_128224448_128224560,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128223720_128223944_128224168,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128223888_128224112_128224056,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128223440_128223608_128223776,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127715424_128223048_128223272,
         output_p1_times_a1_mul_componentxUMxa12_and_b0,
         output_p1_times_a1_mul_componentxUMxcarry_layer2_128223384_128223552,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128223384_128223552,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128222936_128223104_128223216,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128222376_128222600_128222768,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128222432_128222544_128222712,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128221872_128222096_128222264,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128221760_128221928_128222040,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127635584_128221368_128221592,
         output_p1_times_a1_mul_componentxUMxa9_and_b0,
         output_p1_times_a1_mul_componentxUMxsum_layer2_128221424_128221536_128221704,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127827584_127827808_128221256,
         output_p1_times_a1_mul_componentxUMxcarry_layer2_127827752_127827920,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127827752_127827920,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127827248_127827472_127827640,
         output_p1_times_a1_mul_componentxUMxcarry_layer2_127827304_127827416,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127827304_127827416,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127731808_127826912_127827136,
         output_p1_times_a1_mul_componentxUMxa6_and_b0,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127826576_127826800_127826968,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127826464_127826632_127826744,
         output_p1_times_a1_mul_componentxUMxsum_layer2_127672448_127826240_127826520,
         output_p1_times_a1_mul_componentxUMxa3_and_b0,
         output_p1_times_a1_mul_componentxUMxcarry_layer2_127826128_127826296,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127627616_127629520_127824000,
         output_p1_times_a1_mul_componentxUMxa17_and_b0,
         output_p1_times_a1_mul_componentxUMxa16_and_b1,
         output_p1_times_a1_mul_componentxUMxa15_and_b2,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127715984_127849024_127850928,
         output_p1_times_a1_mul_componentxUMxa14_and_b3,
         output_p1_times_a1_mul_componentxUMxa13_and_b4,
         output_p1_times_a1_mul_componentxUMxa12_and_b5,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127636480_127638384_127714080,
         output_p1_times_a1_mul_componentxUMxa11_and_b6,
         output_p1_times_a1_mul_componentxUMxa10_and_b7,
         output_p1_times_a1_mul_componentxUMxa9_and_b8,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127733040_127722720_127724624,
         output_p1_times_a1_mul_componentxUMxa8_and_b9,
         output_p1_times_a1_mul_componentxUMxa7_and_b10,
         output_p1_times_a1_mul_componentxUMxa6_and_b11,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127674016_127675920_127731136,
         output_p1_times_a1_mul_componentxUMxa5_and_b12,
         output_p1_times_a1_mul_componentxUMxa4_and_b13,
         output_p1_times_a1_mul_componentxUMxa3_and_b14,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127832016_127846272_127848176,
         output_p1_times_a1_mul_componentxUMxa2_and_b15,
         output_p1_times_a1_mul_componentxUMxa1_and_b16,
         output_p1_times_a1_mul_componentxUMxa0_and_b17,
         output_p1_times_a1_mul_componentxUMxcarry_layer1_127627504_127629408,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127627504_127629408,
         output_p1_times_a1_mul_componentxUMxa16_and_b0,
         output_p1_times_a1_mul_componentxUMxa15_and_b1,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127715872_127848912_127850816,
         output_p1_times_a1_mul_componentxUMxa14_and_b2,
         output_p1_times_a1_mul_componentxUMxa13_and_b3,
         output_p1_times_a1_mul_componentxUMxa12_and_b4,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127636368_127638272_127713968,
         output_p1_times_a1_mul_componentxUMxa11_and_b5,
         output_p1_times_a1_mul_componentxUMxa10_and_b6,
         output_p1_times_a1_mul_componentxUMxa9_and_b7,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732928_127722608_127724512,
         output_p1_times_a1_mul_componentxUMxa8_and_b8,
         output_p1_times_a1_mul_componentxUMxa7_and_b9,
         output_p1_times_a1_mul_componentxUMxa6_and_b10,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673904_127675808_127731024,
         output_p1_times_a1_mul_componentxUMxa5_and_b11,
         output_p1_times_a1_mul_componentxUMxa4_and_b12,
         output_p1_times_a1_mul_componentxUMxa3_and_b13,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831904_127846160_127848064,
         output_p1_times_a1_mul_componentxUMxa2_and_b14,
         output_p1_times_a1_mul_componentxUMxa1_and_b15,
         output_p1_times_a1_mul_componentxUMxa0_and_b16,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127715760_127848800_127850704,
         output_p1_times_a1_mul_componentxUMxa14_and_b1,
         output_p1_times_a1_mul_componentxUMxa13_and_b2,
         output_p1_times_a1_mul_componentxUMxa12_and_b3,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127636256_127638160_127713856,
         output_p1_times_a1_mul_componentxUMxa11_and_b4,
         output_p1_times_a1_mul_componentxUMxa10_and_b5,
         output_p1_times_a1_mul_componentxUMxa9_and_b6,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732816_127722496_127724400,
         output_p1_times_a1_mul_componentxUMxa8_and_b7,
         output_p1_times_a1_mul_componentxUMxa7_and_b8,
         output_p1_times_a1_mul_componentxUMxa6_and_b9,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673792_127675696_127730912,
         output_p1_times_a1_mul_componentxUMxa5_and_b10,
         output_p1_times_a1_mul_componentxUMxa4_and_b11,
         output_p1_times_a1_mul_componentxUMxa3_and_b12,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831792_127846048_127847952,
         output_p1_times_a1_mul_componentxUMxa2_and_b13,
         output_p1_times_a1_mul_componentxUMxa1_and_b14,
         output_p1_times_a1_mul_componentxUMxa0_and_b15,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127715648_127848688_127850592,
         output_p1_times_a1_mul_componentxUMxa14_and_b0,
         output_p1_times_a1_mul_componentxUMxa13_and_b1,
         output_p1_times_a1_mul_componentxUMxa12_and_b2,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127636144_127638048_127713744,
         output_p1_times_a1_mul_componentxUMxa11_and_b3,
         output_p1_times_a1_mul_componentxUMxa10_and_b4,
         output_p1_times_a1_mul_componentxUMxa9_and_b5,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732704_127722384_127724288,
         output_p1_times_a1_mul_componentxUMxa8_and_b6,
         output_p1_times_a1_mul_componentxUMxa7_and_b7,
         output_p1_times_a1_mul_componentxUMxa6_and_b8,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673680_127675584_127730800,
         output_p1_times_a1_mul_componentxUMxa5_and_b9,
         output_p1_times_a1_mul_componentxUMxa4_and_b10,
         output_p1_times_a1_mul_componentxUMxa3_and_b11,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831680_127845936_127847840,
         output_p1_times_a1_mul_componentxUMxa2_and_b12,
         output_p1_times_a1_mul_componentxUMxa1_and_b13,
         output_p1_times_a1_mul_componentxUMxa0_and_b14,
         output_p1_times_a1_mul_componentxUMxcarry_layer1_127715536_127848576,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127715536_127848576,
         output_p1_times_a1_mul_componentxUMxa13_and_b0,
         output_p1_times_a1_mul_componentxUMxa12_and_b1,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127636032_127637936_127713632,
         output_p1_times_a1_mul_componentxUMxa11_and_b2,
         output_p1_times_a1_mul_componentxUMxa10_and_b3,
         output_p1_times_a1_mul_componentxUMxa9_and_b4,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732592_127722272_127724176,
         output_p1_times_a1_mul_componentxUMxa8_and_b5,
         output_p1_times_a1_mul_componentxUMxa7_and_b6,
         output_p1_times_a1_mul_componentxUMxa6_and_b7,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673568_127675472_127730688,
         output_p1_times_a1_mul_componentxUMxa5_and_b8,
         output_p1_times_a1_mul_componentxUMxa4_and_b9,
         output_p1_times_a1_mul_componentxUMxa3_and_b10,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831568_127845824_127847728,
         output_p1_times_a1_mul_componentxUMxa2_and_b11,
         output_p1_times_a1_mul_componentxUMxa1_and_b12,
         output_p1_times_a1_mul_componentxUMxa0_and_b13,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127635920_127637824_127713520,
         output_p1_times_a1_mul_componentxUMxa11_and_b1,
         output_p1_times_a1_mul_componentxUMxa10_and_b2,
         output_p1_times_a1_mul_componentxUMxa9_and_b3,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732480_127722160_127724064,
         output_p1_times_a1_mul_componentxUMxa8_and_b4,
         output_p1_times_a1_mul_componentxUMxa7_and_b5,
         output_p1_times_a1_mul_componentxUMxa6_and_b6,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673456_127675360_127730576,
         output_p1_times_a1_mul_componentxUMxa5_and_b7,
         output_p1_times_a1_mul_componentxUMxa4_and_b8,
         output_p1_times_a1_mul_componentxUMxa3_and_b9,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831456_127845712_127847616,
         output_p1_times_a1_mul_componentxUMxa2_and_b10,
         output_p1_times_a1_mul_componentxUMxa1_and_b11,
         output_p1_times_a1_mul_componentxUMxa0_and_b12,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127635808_127637712_127713408,
         output_p1_times_a1_mul_componentxUMxa11_and_b0,
         output_p1_times_a1_mul_componentxUMxa10_and_b1,
         output_p1_times_a1_mul_componentxUMxa9_and_b2,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732368_127722048_127723952,
         output_p1_times_a1_mul_componentxUMxa8_and_b3,
         output_p1_times_a1_mul_componentxUMxa7_and_b4,
         output_p1_times_a1_mul_componentxUMxa6_and_b5,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673344_127675248_127730464,
         output_p1_times_a1_mul_componentxUMxa5_and_b6,
         output_p1_times_a1_mul_componentxUMxa4_and_b7,
         output_p1_times_a1_mul_componentxUMxa3_and_b8,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831344_127845600_127847504,
         output_p1_times_a1_mul_componentxUMxa2_and_b9,
         output_p1_times_a1_mul_componentxUMxa1_and_b10,
         output_p1_times_a1_mul_componentxUMxa0_and_b11,
         output_p1_times_a1_mul_componentxUMxcarry_layer1_127635696_127637600,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127635696_127637600,
         output_p1_times_a1_mul_componentxUMxa10_and_b0,
         output_p1_times_a1_mul_componentxUMxa9_and_b1,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732256_127721936_127723840,
         output_p1_times_a1_mul_componentxUMxa8_and_b2,
         output_p1_times_a1_mul_componentxUMxa7_and_b3,
         output_p1_times_a1_mul_componentxUMxa6_and_b4,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673232_127675136_127730352,
         output_p1_times_a1_mul_componentxUMxa5_and_b5,
         output_p1_times_a1_mul_componentxUMxa4_and_b6,
         output_p1_times_a1_mul_componentxUMxa3_and_b7,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831232_127845488_127847392,
         output_p1_times_a1_mul_componentxUMxa2_and_b8,
         output_p1_times_a1_mul_componentxUMxa1_and_b9,
         output_p1_times_a1_mul_componentxUMxa0_and_b10,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732144_127721824_127723728,
         output_p1_times_a1_mul_componentxUMxa8_and_b1,
         output_p1_times_a1_mul_componentxUMxa7_and_b2,
         output_p1_times_a1_mul_componentxUMxa6_and_b3,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673120_127675024_127730240,
         output_p1_times_a1_mul_componentxUMxa5_and_b4,
         output_p1_times_a1_mul_componentxUMxa4_and_b5,
         output_p1_times_a1_mul_componentxUMxa3_and_b6,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831120_127845376_127847280,
         output_p1_times_a1_mul_componentxUMxa2_and_b7,
         output_p1_times_a1_mul_componentxUMxa1_and_b8,
         output_p1_times_a1_mul_componentxUMxa0_and_b9,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127732032_127721712_127723616,
         output_p1_times_a1_mul_componentxUMxa8_and_b0,
         output_p1_times_a1_mul_componentxUMxa7_and_b1,
         output_p1_times_a1_mul_componentxUMxa6_and_b2,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127673008_127674912_127730128,
         output_p1_times_a1_mul_componentxUMxa5_and_b3,
         output_p1_times_a1_mul_componentxUMxa4_and_b4,
         output_p1_times_a1_mul_componentxUMxa3_and_b5,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127831008_127845264_127847168,
         output_p1_times_a1_mul_componentxUMxa2_and_b6,
         output_p1_times_a1_mul_componentxUMxa1_and_b7,
         output_p1_times_a1_mul_componentxUMxa0_and_b8,
         output_p1_times_a1_mul_componentxUMxcarry_layer1_127731920_127721600,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127731920_127721600,
         output_p1_times_a1_mul_componentxUMxa7_and_b0,
         output_p1_times_a1_mul_componentxUMxa6_and_b1,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127672896_127674800_127730016,
         output_p1_times_a1_mul_componentxUMxa5_and_b2,
         output_p1_times_a1_mul_componentxUMxa4_and_b3,
         output_p1_times_a1_mul_componentxUMxa3_and_b4,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127830896_127845152_127847056,
         output_p1_times_a1_mul_componentxUMxa2_and_b5,
         output_p1_times_a1_mul_componentxUMxa1_and_b6,
         output_p1_times_a1_mul_componentxUMxa0_and_b7,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127672784_127674688_127729904,
         output_p1_times_a1_mul_componentxUMxa5_and_b1,
         output_p1_times_a1_mul_componentxUMxa4_and_b2,
         output_p1_times_a1_mul_componentxUMxa3_and_b3,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127830784_127845040_127846944,
         output_p1_times_a1_mul_componentxUMxa2_and_b4,
         output_p1_times_a1_mul_componentxUMxa1_and_b5,
         output_p1_times_a1_mul_componentxUMxa0_and_b6,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127672672_127674576_127729792,
         output_p1_times_a1_mul_componentxUMxa5_and_b0,
         output_p1_times_a1_mul_componentxUMxa4_and_b1,
         output_p1_times_a1_mul_componentxUMxa3_and_b2,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127830672_127844928_127846832,
         output_p1_times_a1_mul_componentxUMxa2_and_b3,
         output_p1_times_a1_mul_componentxUMxa1_and_b4,
         output_p1_times_a1_mul_componentxUMxa0_and_b5,
         output_p1_times_a1_mul_componentxUMxcarry_layer1_127672560_127674464,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127672560_127674464,
         output_p1_times_a1_mul_componentxUMxa4_and_b0,
         output_p1_times_a1_mul_componentxUMxa3_and_b1,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127830560_127844816_127846720,
         output_p1_times_a1_mul_componentxUMxa2_and_b2,
         output_p1_times_a1_mul_componentxUMxa1_and_b3,
         output_p1_times_a1_mul_componentxUMxa0_and_b4,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127830448_127844704_127846608,
         output_p1_times_a1_mul_componentxUMxa2_and_b1,
         output_p1_times_a1_mul_componentxUMxa1_and_b2,
         output_p1_times_a1_mul_componentxUMxa0_and_b3,
         output_p1_times_a1_mul_componentxUMxsum_layer1_127830336_127844592_127846496,
         output_p1_times_a1_mul_componentxUMxa2_and_b0,
         output_p1_times_a1_mul_componentxUMxa1_and_b1,
         output_p1_times_a1_mul_componentxUMxa0_and_b2,
         output_p1_times_a1_mul_componentxUMxcarry_layer1_127830168_127844480,
         output_p1_times_a1_mul_componentxUMxa1_and_b0,
         output_p1_times_a1_mul_componentxUMxa0_and_b1,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128315744_128315968_128316136,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128315464_128315632_128315800,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128220800_128221024_128221136,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128220688_128220856_128220968,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128126256_128220520_128220744,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128125920_128220352_128220576,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128125584_128220184_128220408,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128125248_128219960_128220240,
         input_p2_times_b2_mul_componentxUMxcarry_layer5_128219792_128220016,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128219792_128220016,
         input_p2_times_b2_mul_componentxUMxcarry_layer5_128219624_128219848,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128219624_128219848,
         input_p2_times_b2_mul_componentxUMxcarry_layer5_128219456_128219680,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128219456_128219680,
         input_p2_times_b2_mul_componentxUMxcarry_layer5_128219288_128219512,
         input_p2_times_b2_mul_componentxUMxsum_layer5_128219288_128219512,
         input_p2_times_b2_mul_componentxUMxcarry_layer5_128219120_128219344,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128238312_128238424_128238592,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128237752_128237976_128238144,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128237920_128238088,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128126760_128237640_128237808,
         input_p2_times_b2_mul_componentxUMxcarry_layer4_128126816_128126928,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128126816_128126928,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128263168_128126424_128126648,
         input_p2_times_b2_mul_componentxUMxcarry_layer4_128126480_128126592,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128126480_128126592,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128262496_128126088_128126312,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128125752_128125976_128126144,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128125416_128125640_128125808,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128125080_128125304_128125472,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128124744_128124968_128125136,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128124632_128124800_128124912,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128247456_128124464_128124688,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128247120_128124240_128124520,
         input_p2_times_b2_mul_componentxUMxcarry_layer4_128124072_128124296,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128124072_128124296,
         input_p2_times_b2_mul_componentxUMxcarry_layer4_128123904_128124128,
         input_p2_times_b2_mul_componentxUMxsum_layer4_128123904_128124128,
         input_p2_times_b2_mul_componentxUMxcarry_layer4_128123792_128123960,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128264344_128264512,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128263896_128264064_128264176,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128263336_128263560_128263728,
         input_p2_times_b2_mul_componentxUMxcarry_layer3_128263672_128263840,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128263672_128263840,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128263224_128263392_128263504,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128262664_128262888_128263056,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128262720_128262832_128263000,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128262216_128262384_128262552,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128249696_128249808_128262328,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128197128_128249304_128249528,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128249360_128249472_128249640,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128248800_128249024_128249192,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128248856_128248968_128249136,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128248296_128248520_128248688,
         input_p2_times_b2_mul_componentxUMxcarry_layer3_128248464_128248632,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128248464_128248632,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128247960_128248184_128248352,
         input_p2_times_b2_mul_componentxUMxcarry_layer3_128248016_128248128,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128248016_128248128,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128222880_128247624_128247848,
         input_p2_times_b2_mul_componentxUMxcarry_layer3_128247680_128247792,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128247680_128247792,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128222208_128247288_128247512,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128246952_128247176_128247344,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128246616_128246840_128247008,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128246504_128246672_128246784,
         input_p2_times_b2_mul_componentxUMxsum_layer3_127827080_128246280_128246560,
         input_p2_times_b2_mul_componentxUMxcarry_layer3_128246112_128246336,
         input_p2_times_b2_mul_componentxUMxsum_layer3_128246112_128246336,
         input_p2_times_b2_mul_componentxUMxcarry_layer3_128246000_128246168,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128199816_128200040_128199984,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128199368_128199480_128199648,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128198864_128199032_128199200,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128198304_128198528_128198696,
         input_p2_times_b2_mul_componentxUMxcarry_layer2_128198976_128199144,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128198976_128199144,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128198472_128198640_128198808,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128198080_128198192_128198360,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128197464_128197688_128197856,
         input_p2_times_b2_mul_componentxUMxcarry_layer2_128198024_128197968,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128198024_128197968,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128197520_128197632_128197800,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128197016_128197240_128197352,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127627392_128196680_128196848,
         input_p2_times_b2_mul_componentxUMxa15_and_b0,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128196792_128196960_128197184,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128224952_128225120_128225232,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128224392_128224616_128224784,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128224728_128224896_128225064,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128224280_128224448_128224560,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128223720_128223944_128224168,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128223888_128224112_128224056,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128223440_128223608_128223776,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127715424_128223048_128223272,
         input_p2_times_b2_mul_componentxUMxa12_and_b0,
         input_p2_times_b2_mul_componentxUMxcarry_layer2_128223384_128223552,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128223384_128223552,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128222936_128223104_128223216,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128222376_128222600_128222768,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128222432_128222544_128222712,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128221872_128222096_128222264,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128221760_128221928_128222040,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127635584_128221368_128221592,
         input_p2_times_b2_mul_componentxUMxa9_and_b0,
         input_p2_times_b2_mul_componentxUMxsum_layer2_128221424_128221536_128221704,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127827584_127827808_128221256,
         input_p2_times_b2_mul_componentxUMxcarry_layer2_127827752_127827920,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127827752_127827920,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127827248_127827472_127827640,
         input_p2_times_b2_mul_componentxUMxcarry_layer2_127827304_127827416,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127827304_127827416,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127731808_127826912_127827136,
         input_p2_times_b2_mul_componentxUMxa6_and_b0,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127826576_127826800_127826968,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127826464_127826632_127826744,
         input_p2_times_b2_mul_componentxUMxsum_layer2_127672448_127826240_127826520,
         input_p2_times_b2_mul_componentxUMxa3_and_b0,
         input_p2_times_b2_mul_componentxUMxcarry_layer2_127826128_127826296,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127627616_127629520_127824000,
         input_p2_times_b2_mul_componentxUMxa17_and_b0,
         input_p2_times_b2_mul_componentxUMxa16_and_b1,
         input_p2_times_b2_mul_componentxUMxa15_and_b2,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127715984_127849024_127850928,
         input_p2_times_b2_mul_componentxUMxa14_and_b3,
         input_p2_times_b2_mul_componentxUMxa13_and_b4,
         input_p2_times_b2_mul_componentxUMxa12_and_b5,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127636480_127638384_127714080,
         input_p2_times_b2_mul_componentxUMxa11_and_b6,
         input_p2_times_b2_mul_componentxUMxa10_and_b7,
         input_p2_times_b2_mul_componentxUMxa9_and_b8,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127733040_127722720_127724624,
         input_p2_times_b2_mul_componentxUMxa8_and_b9,
         input_p2_times_b2_mul_componentxUMxa7_and_b10,
         input_p2_times_b2_mul_componentxUMxa6_and_b11,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127674016_127675920_127731136,
         input_p2_times_b2_mul_componentxUMxa5_and_b12,
         input_p2_times_b2_mul_componentxUMxa4_and_b13,
         input_p2_times_b2_mul_componentxUMxa3_and_b14,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127832016_127846272_127848176,
         input_p2_times_b2_mul_componentxUMxa2_and_b15,
         input_p2_times_b2_mul_componentxUMxa1_and_b16,
         input_p2_times_b2_mul_componentxUMxa0_and_b17,
         input_p2_times_b2_mul_componentxUMxcarry_layer1_127627504_127629408,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127627504_127629408,
         input_p2_times_b2_mul_componentxUMxa16_and_b0,
         input_p2_times_b2_mul_componentxUMxa15_and_b1,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127715872_127848912_127850816,
         input_p2_times_b2_mul_componentxUMxa14_and_b2,
         input_p2_times_b2_mul_componentxUMxa13_and_b3,
         input_p2_times_b2_mul_componentxUMxa12_and_b4,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127636368_127638272_127713968,
         input_p2_times_b2_mul_componentxUMxa11_and_b5,
         input_p2_times_b2_mul_componentxUMxa10_and_b6,
         input_p2_times_b2_mul_componentxUMxa9_and_b7,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732928_127722608_127724512,
         input_p2_times_b2_mul_componentxUMxa8_and_b8,
         input_p2_times_b2_mul_componentxUMxa7_and_b9,
         input_p2_times_b2_mul_componentxUMxa6_and_b10,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673904_127675808_127731024,
         input_p2_times_b2_mul_componentxUMxa5_and_b11,
         input_p2_times_b2_mul_componentxUMxa4_and_b12,
         input_p2_times_b2_mul_componentxUMxa3_and_b13,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831904_127846160_127848064,
         input_p2_times_b2_mul_componentxUMxa2_and_b14,
         input_p2_times_b2_mul_componentxUMxa1_and_b15,
         input_p2_times_b2_mul_componentxUMxa0_and_b16,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127715760_127848800_127850704,
         input_p2_times_b2_mul_componentxUMxa14_and_b1,
         input_p2_times_b2_mul_componentxUMxa13_and_b2,
         input_p2_times_b2_mul_componentxUMxa12_and_b3,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127636256_127638160_127713856,
         input_p2_times_b2_mul_componentxUMxa11_and_b4,
         input_p2_times_b2_mul_componentxUMxa10_and_b5,
         input_p2_times_b2_mul_componentxUMxa9_and_b6,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732816_127722496_127724400,
         input_p2_times_b2_mul_componentxUMxa8_and_b7,
         input_p2_times_b2_mul_componentxUMxa7_and_b8,
         input_p2_times_b2_mul_componentxUMxa6_and_b9,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673792_127675696_127730912,
         input_p2_times_b2_mul_componentxUMxa5_and_b10,
         input_p2_times_b2_mul_componentxUMxa4_and_b11,
         input_p2_times_b2_mul_componentxUMxa3_and_b12,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831792_127846048_127847952,
         input_p2_times_b2_mul_componentxUMxa2_and_b13,
         input_p2_times_b2_mul_componentxUMxa1_and_b14,
         input_p2_times_b2_mul_componentxUMxa0_and_b15,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127715648_127848688_127850592,
         input_p2_times_b2_mul_componentxUMxa14_and_b0,
         input_p2_times_b2_mul_componentxUMxa13_and_b1,
         input_p2_times_b2_mul_componentxUMxa12_and_b2,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127636144_127638048_127713744,
         input_p2_times_b2_mul_componentxUMxa11_and_b3,
         input_p2_times_b2_mul_componentxUMxa10_and_b4,
         input_p2_times_b2_mul_componentxUMxa9_and_b5,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732704_127722384_127724288,
         input_p2_times_b2_mul_componentxUMxa8_and_b6,
         input_p2_times_b2_mul_componentxUMxa7_and_b7,
         input_p2_times_b2_mul_componentxUMxa6_and_b8,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673680_127675584_127730800,
         input_p2_times_b2_mul_componentxUMxa5_and_b9,
         input_p2_times_b2_mul_componentxUMxa4_and_b10,
         input_p2_times_b2_mul_componentxUMxa3_and_b11,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831680_127845936_127847840,
         input_p2_times_b2_mul_componentxUMxa2_and_b12,
         input_p2_times_b2_mul_componentxUMxa1_and_b13,
         input_p2_times_b2_mul_componentxUMxa0_and_b14,
         input_p2_times_b2_mul_componentxUMxcarry_layer1_127715536_127848576,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127715536_127848576,
         input_p2_times_b2_mul_componentxUMxa13_and_b0,
         input_p2_times_b2_mul_componentxUMxa12_and_b1,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127636032_127637936_127713632,
         input_p2_times_b2_mul_componentxUMxa11_and_b2,
         input_p2_times_b2_mul_componentxUMxa10_and_b3,
         input_p2_times_b2_mul_componentxUMxa9_and_b4,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732592_127722272_127724176,
         input_p2_times_b2_mul_componentxUMxa8_and_b5,
         input_p2_times_b2_mul_componentxUMxa7_and_b6,
         input_p2_times_b2_mul_componentxUMxa6_and_b7,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673568_127675472_127730688,
         input_p2_times_b2_mul_componentxUMxa5_and_b8,
         input_p2_times_b2_mul_componentxUMxa4_and_b9,
         input_p2_times_b2_mul_componentxUMxa3_and_b10,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831568_127845824_127847728,
         input_p2_times_b2_mul_componentxUMxa2_and_b11,
         input_p2_times_b2_mul_componentxUMxa1_and_b12,
         input_p2_times_b2_mul_componentxUMxa0_and_b13,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127635920_127637824_127713520,
         input_p2_times_b2_mul_componentxUMxa11_and_b1,
         input_p2_times_b2_mul_componentxUMxa10_and_b2,
         input_p2_times_b2_mul_componentxUMxa9_and_b3,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732480_127722160_127724064,
         input_p2_times_b2_mul_componentxUMxa8_and_b4,
         input_p2_times_b2_mul_componentxUMxa7_and_b5,
         input_p2_times_b2_mul_componentxUMxa6_and_b6,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673456_127675360_127730576,
         input_p2_times_b2_mul_componentxUMxa5_and_b7,
         input_p2_times_b2_mul_componentxUMxa4_and_b8,
         input_p2_times_b2_mul_componentxUMxa3_and_b9,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831456_127845712_127847616,
         input_p2_times_b2_mul_componentxUMxa2_and_b10,
         input_p2_times_b2_mul_componentxUMxa1_and_b11,
         input_p2_times_b2_mul_componentxUMxa0_and_b12,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127635808_127637712_127713408,
         input_p2_times_b2_mul_componentxUMxa11_and_b0,
         input_p2_times_b2_mul_componentxUMxa10_and_b1,
         input_p2_times_b2_mul_componentxUMxa9_and_b2,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732368_127722048_127723952,
         input_p2_times_b2_mul_componentxUMxa8_and_b3,
         input_p2_times_b2_mul_componentxUMxa7_and_b4,
         input_p2_times_b2_mul_componentxUMxa6_and_b5,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673344_127675248_127730464,
         input_p2_times_b2_mul_componentxUMxa5_and_b6,
         input_p2_times_b2_mul_componentxUMxa4_and_b7,
         input_p2_times_b2_mul_componentxUMxa3_and_b8,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831344_127845600_127847504,
         input_p2_times_b2_mul_componentxUMxa2_and_b9,
         input_p2_times_b2_mul_componentxUMxa1_and_b10,
         input_p2_times_b2_mul_componentxUMxa0_and_b11,
         input_p2_times_b2_mul_componentxUMxcarry_layer1_127635696_127637600,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127635696_127637600,
         input_p2_times_b2_mul_componentxUMxa10_and_b0,
         input_p2_times_b2_mul_componentxUMxa9_and_b1,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732256_127721936_127723840,
         input_p2_times_b2_mul_componentxUMxa8_and_b2,
         input_p2_times_b2_mul_componentxUMxa7_and_b3,
         input_p2_times_b2_mul_componentxUMxa6_and_b4,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673232_127675136_127730352,
         input_p2_times_b2_mul_componentxUMxa5_and_b5,
         input_p2_times_b2_mul_componentxUMxa4_and_b6,
         input_p2_times_b2_mul_componentxUMxa3_and_b7,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831232_127845488_127847392,
         input_p2_times_b2_mul_componentxUMxa2_and_b8,
         input_p2_times_b2_mul_componentxUMxa1_and_b9,
         input_p2_times_b2_mul_componentxUMxa0_and_b10,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732144_127721824_127723728,
         input_p2_times_b2_mul_componentxUMxa8_and_b1,
         input_p2_times_b2_mul_componentxUMxa7_and_b2,
         input_p2_times_b2_mul_componentxUMxa6_and_b3,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673120_127675024_127730240,
         input_p2_times_b2_mul_componentxUMxa5_and_b4,
         input_p2_times_b2_mul_componentxUMxa4_and_b5,
         input_p2_times_b2_mul_componentxUMxa3_and_b6,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831120_127845376_127847280,
         input_p2_times_b2_mul_componentxUMxa2_and_b7,
         input_p2_times_b2_mul_componentxUMxa1_and_b8,
         input_p2_times_b2_mul_componentxUMxa0_and_b9,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127732032_127721712_127723616,
         input_p2_times_b2_mul_componentxUMxa8_and_b0,
         input_p2_times_b2_mul_componentxUMxa7_and_b1,
         input_p2_times_b2_mul_componentxUMxa6_and_b2,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127673008_127674912_127730128,
         input_p2_times_b2_mul_componentxUMxa5_and_b3,
         input_p2_times_b2_mul_componentxUMxa4_and_b4,
         input_p2_times_b2_mul_componentxUMxa3_and_b5,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127831008_127845264_127847168,
         input_p2_times_b2_mul_componentxUMxa2_and_b6,
         input_p2_times_b2_mul_componentxUMxa1_and_b7,
         input_p2_times_b2_mul_componentxUMxa0_and_b8,
         input_p2_times_b2_mul_componentxUMxcarry_layer1_127731920_127721600,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127731920_127721600,
         input_p2_times_b2_mul_componentxUMxa7_and_b0,
         input_p2_times_b2_mul_componentxUMxa6_and_b1,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127672896_127674800_127730016,
         input_p2_times_b2_mul_componentxUMxa5_and_b2,
         input_p2_times_b2_mul_componentxUMxa4_and_b3,
         input_p2_times_b2_mul_componentxUMxa3_and_b4,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127830896_127845152_127847056,
         input_p2_times_b2_mul_componentxUMxa2_and_b5,
         input_p2_times_b2_mul_componentxUMxa1_and_b6,
         input_p2_times_b2_mul_componentxUMxa0_and_b7,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127672784_127674688_127729904,
         input_p2_times_b2_mul_componentxUMxa5_and_b1,
         input_p2_times_b2_mul_componentxUMxa4_and_b2,
         input_p2_times_b2_mul_componentxUMxa3_and_b3,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127830784_127845040_127846944,
         input_p2_times_b2_mul_componentxUMxa2_and_b4,
         input_p2_times_b2_mul_componentxUMxa1_and_b5,
         input_p2_times_b2_mul_componentxUMxa0_and_b6,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127672672_127674576_127729792,
         input_p2_times_b2_mul_componentxUMxa5_and_b0,
         input_p2_times_b2_mul_componentxUMxa4_and_b1,
         input_p2_times_b2_mul_componentxUMxa3_and_b2,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127830672_127844928_127846832,
         input_p2_times_b2_mul_componentxUMxa2_and_b3,
         input_p2_times_b2_mul_componentxUMxa1_and_b4,
         input_p2_times_b2_mul_componentxUMxa0_and_b5,
         input_p2_times_b2_mul_componentxUMxcarry_layer1_127672560_127674464,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127672560_127674464,
         input_p2_times_b2_mul_componentxUMxa4_and_b0,
         input_p2_times_b2_mul_componentxUMxa3_and_b1,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127830560_127844816_127846720,
         input_p2_times_b2_mul_componentxUMxa2_and_b2,
         input_p2_times_b2_mul_componentxUMxa1_and_b3,
         input_p2_times_b2_mul_componentxUMxa0_and_b4,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127830448_127844704_127846608,
         input_p2_times_b2_mul_componentxUMxa2_and_b1,
         input_p2_times_b2_mul_componentxUMxa1_and_b2,
         input_p2_times_b2_mul_componentxUMxa0_and_b3,
         input_p2_times_b2_mul_componentxUMxsum_layer1_127830336_127844592_127846496,
         input_p2_times_b2_mul_componentxUMxa2_and_b0,
         input_p2_times_b2_mul_componentxUMxa1_and_b1,
         input_p2_times_b2_mul_componentxUMxa0_and_b2,
         input_p2_times_b2_mul_componentxUMxcarry_layer1_127830168_127844480,
         input_p2_times_b2_mul_componentxUMxa1_and_b0,
         input_p2_times_b2_mul_componentxUMxa0_and_b1,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128315744_128315968_128316136,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128315464_128315632_128315800,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128220800_128221024_128221136,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128220688_128220856_128220968,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128126256_128220520_128220744,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128125920_128220352_128220576,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128125584_128220184_128220408,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128125248_128219960_128220240,
         input_p1_times_b1_mul_componentxUMxcarry_layer5_128219792_128220016,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128219792_128220016,
         input_p1_times_b1_mul_componentxUMxcarry_layer5_128219624_128219848,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128219624_128219848,
         input_p1_times_b1_mul_componentxUMxcarry_layer5_128219456_128219680,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128219456_128219680,
         input_p1_times_b1_mul_componentxUMxcarry_layer5_128219288_128219512,
         input_p1_times_b1_mul_componentxUMxsum_layer5_128219288_128219512,
         input_p1_times_b1_mul_componentxUMxcarry_layer5_128219120_128219344,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128238312_128238424_128238592,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128237752_128237976_128238144,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128237920_128238088,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128126760_128237640_128237808,
         input_p1_times_b1_mul_componentxUMxcarry_layer4_128126816_128126928,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128126816_128126928,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128263168_128126424_128126648,
         input_p1_times_b1_mul_componentxUMxcarry_layer4_128126480_128126592,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128126480_128126592,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128262496_128126088_128126312,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128125752_128125976_128126144,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128125416_128125640_128125808,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128125080_128125304_128125472,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128124744_128124968_128125136,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128124632_128124800_128124912,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128247456_128124464_128124688,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128247120_128124240_128124520,
         input_p1_times_b1_mul_componentxUMxcarry_layer4_128124072_128124296,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128124072_128124296,
         input_p1_times_b1_mul_componentxUMxcarry_layer4_128123904_128124128,
         input_p1_times_b1_mul_componentxUMxsum_layer4_128123904_128124128,
         input_p1_times_b1_mul_componentxUMxcarry_layer4_128123792_128123960,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128264344_128264512,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128263896_128264064_128264176,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128263336_128263560_128263728,
         input_p1_times_b1_mul_componentxUMxcarry_layer3_128263672_128263840,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128263672_128263840,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128263224_128263392_128263504,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128262664_128262888_128263056,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128262720_128262832_128263000,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128262216_128262384_128262552,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128249696_128249808_128262328,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128197128_128249304_128249528,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128249360_128249472_128249640,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128248800_128249024_128249192,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128248856_128248968_128249136,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128248296_128248520_128248688,
         input_p1_times_b1_mul_componentxUMxcarry_layer3_128248464_128248632,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128248464_128248632,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128247960_128248184_128248352,
         input_p1_times_b1_mul_componentxUMxcarry_layer3_128248016_128248128,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128248016_128248128,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128222880_128247624_128247848,
         input_p1_times_b1_mul_componentxUMxcarry_layer3_128247680_128247792,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128247680_128247792,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128222208_128247288_128247512,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128246952_128247176_128247344,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128246616_128246840_128247008,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128246504_128246672_128246784,
         input_p1_times_b1_mul_componentxUMxsum_layer3_127827080_128246280_128246560,
         input_p1_times_b1_mul_componentxUMxcarry_layer3_128246112_128246336,
         input_p1_times_b1_mul_componentxUMxsum_layer3_128246112_128246336,
         input_p1_times_b1_mul_componentxUMxcarry_layer3_128246000_128246168,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128199816_128200040_128199984,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128199368_128199480_128199648,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128198864_128199032_128199200,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128198304_128198528_128198696,
         input_p1_times_b1_mul_componentxUMxcarry_layer2_128198976_128199144,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128198976_128199144,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128198472_128198640_128198808,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128198080_128198192_128198360,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128197464_128197688_128197856,
         input_p1_times_b1_mul_componentxUMxcarry_layer2_128198024_128197968,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128198024_128197968,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128197520_128197632_128197800,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128197016_128197240_128197352,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127627392_128196680_128196848,
         input_p1_times_b1_mul_componentxUMxa15_and_b0,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128196792_128196960_128197184,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128224952_128225120_128225232,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128224392_128224616_128224784,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128224728_128224896_128225064,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128224280_128224448_128224560,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128223720_128223944_128224168,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128223888_128224112_128224056,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128223440_128223608_128223776,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127715424_128223048_128223272,
         input_p1_times_b1_mul_componentxUMxa12_and_b0,
         input_p1_times_b1_mul_componentxUMxcarry_layer2_128223384_128223552,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128223384_128223552,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128222936_128223104_128223216,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128222376_128222600_128222768,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128222432_128222544_128222712,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128221872_128222096_128222264,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128221760_128221928_128222040,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127635584_128221368_128221592,
         input_p1_times_b1_mul_componentxUMxa9_and_b0,
         input_p1_times_b1_mul_componentxUMxsum_layer2_128221424_128221536_128221704,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127827584_127827808_128221256,
         input_p1_times_b1_mul_componentxUMxcarry_layer2_127827752_127827920,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127827752_127827920,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127827248_127827472_127827640,
         input_p1_times_b1_mul_componentxUMxcarry_layer2_127827304_127827416,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127827304_127827416,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127731808_127826912_127827136,
         input_p1_times_b1_mul_componentxUMxa6_and_b0,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127826576_127826800_127826968,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127826464_127826632_127826744,
         input_p1_times_b1_mul_componentxUMxsum_layer2_127672448_127826240_127826520,
         input_p1_times_b1_mul_componentxUMxa3_and_b0,
         input_p1_times_b1_mul_componentxUMxcarry_layer2_127826128_127826296,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127627616_127629520_127824000,
         input_p1_times_b1_mul_componentxUMxa17_and_b0,
         input_p1_times_b1_mul_componentxUMxa16_and_b1,
         input_p1_times_b1_mul_componentxUMxa15_and_b2,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127715984_127849024_127850928,
         input_p1_times_b1_mul_componentxUMxa14_and_b3,
         input_p1_times_b1_mul_componentxUMxa13_and_b4,
         input_p1_times_b1_mul_componentxUMxa12_and_b5,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127636480_127638384_127714080,
         input_p1_times_b1_mul_componentxUMxa11_and_b6,
         input_p1_times_b1_mul_componentxUMxa10_and_b7,
         input_p1_times_b1_mul_componentxUMxa9_and_b8,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127733040_127722720_127724624,
         input_p1_times_b1_mul_componentxUMxa8_and_b9,
         input_p1_times_b1_mul_componentxUMxa7_and_b10,
         input_p1_times_b1_mul_componentxUMxa6_and_b11,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127674016_127675920_127731136,
         input_p1_times_b1_mul_componentxUMxa5_and_b12,
         input_p1_times_b1_mul_componentxUMxa4_and_b13,
         input_p1_times_b1_mul_componentxUMxa3_and_b14,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127832016_127846272_127848176,
         input_p1_times_b1_mul_componentxUMxa2_and_b15,
         input_p1_times_b1_mul_componentxUMxa1_and_b16,
         input_p1_times_b1_mul_componentxUMxa0_and_b17,
         input_p1_times_b1_mul_componentxUMxcarry_layer1_127627504_127629408,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127627504_127629408,
         input_p1_times_b1_mul_componentxUMxa16_and_b0,
         input_p1_times_b1_mul_componentxUMxa15_and_b1,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127715872_127848912_127850816,
         input_p1_times_b1_mul_componentxUMxa14_and_b2,
         input_p1_times_b1_mul_componentxUMxa13_and_b3,
         input_p1_times_b1_mul_componentxUMxa12_and_b4,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127636368_127638272_127713968,
         input_p1_times_b1_mul_componentxUMxa11_and_b5,
         input_p1_times_b1_mul_componentxUMxa10_and_b6,
         input_p1_times_b1_mul_componentxUMxa9_and_b7,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732928_127722608_127724512,
         input_p1_times_b1_mul_componentxUMxa8_and_b8,
         input_p1_times_b1_mul_componentxUMxa7_and_b9,
         input_p1_times_b1_mul_componentxUMxa6_and_b10,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673904_127675808_127731024,
         input_p1_times_b1_mul_componentxUMxa5_and_b11,
         input_p1_times_b1_mul_componentxUMxa4_and_b12,
         input_p1_times_b1_mul_componentxUMxa3_and_b13,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831904_127846160_127848064,
         input_p1_times_b1_mul_componentxUMxa2_and_b14,
         input_p1_times_b1_mul_componentxUMxa1_and_b15,
         input_p1_times_b1_mul_componentxUMxa0_and_b16,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127715760_127848800_127850704,
         input_p1_times_b1_mul_componentxUMxa14_and_b1,
         input_p1_times_b1_mul_componentxUMxa13_and_b2,
         input_p1_times_b1_mul_componentxUMxa12_and_b3,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127636256_127638160_127713856,
         input_p1_times_b1_mul_componentxUMxa11_and_b4,
         input_p1_times_b1_mul_componentxUMxa10_and_b5,
         input_p1_times_b1_mul_componentxUMxa9_and_b6,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732816_127722496_127724400,
         input_p1_times_b1_mul_componentxUMxa8_and_b7,
         input_p1_times_b1_mul_componentxUMxa7_and_b8,
         input_p1_times_b1_mul_componentxUMxa6_and_b9,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673792_127675696_127730912,
         input_p1_times_b1_mul_componentxUMxa5_and_b10,
         input_p1_times_b1_mul_componentxUMxa4_and_b11,
         input_p1_times_b1_mul_componentxUMxa3_and_b12,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831792_127846048_127847952,
         input_p1_times_b1_mul_componentxUMxa2_and_b13,
         input_p1_times_b1_mul_componentxUMxa1_and_b14,
         input_p1_times_b1_mul_componentxUMxa0_and_b15,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127715648_127848688_127850592,
         input_p1_times_b1_mul_componentxUMxa14_and_b0,
         input_p1_times_b1_mul_componentxUMxa13_and_b1,
         input_p1_times_b1_mul_componentxUMxa12_and_b2,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127636144_127638048_127713744,
         input_p1_times_b1_mul_componentxUMxa11_and_b3,
         input_p1_times_b1_mul_componentxUMxa10_and_b4,
         input_p1_times_b1_mul_componentxUMxa9_and_b5,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732704_127722384_127724288,
         input_p1_times_b1_mul_componentxUMxa8_and_b6,
         input_p1_times_b1_mul_componentxUMxa7_and_b7,
         input_p1_times_b1_mul_componentxUMxa6_and_b8,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673680_127675584_127730800,
         input_p1_times_b1_mul_componentxUMxa5_and_b9,
         input_p1_times_b1_mul_componentxUMxa4_and_b10,
         input_p1_times_b1_mul_componentxUMxa3_and_b11,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831680_127845936_127847840,
         input_p1_times_b1_mul_componentxUMxa2_and_b12,
         input_p1_times_b1_mul_componentxUMxa1_and_b13,
         input_p1_times_b1_mul_componentxUMxa0_and_b14,
         input_p1_times_b1_mul_componentxUMxcarry_layer1_127715536_127848576,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127715536_127848576,
         input_p1_times_b1_mul_componentxUMxa13_and_b0,
         input_p1_times_b1_mul_componentxUMxa12_and_b1,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127636032_127637936_127713632,
         input_p1_times_b1_mul_componentxUMxa11_and_b2,
         input_p1_times_b1_mul_componentxUMxa10_and_b3,
         input_p1_times_b1_mul_componentxUMxa9_and_b4,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732592_127722272_127724176,
         input_p1_times_b1_mul_componentxUMxa8_and_b5,
         input_p1_times_b1_mul_componentxUMxa7_and_b6,
         input_p1_times_b1_mul_componentxUMxa6_and_b7,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673568_127675472_127730688,
         input_p1_times_b1_mul_componentxUMxa5_and_b8,
         input_p1_times_b1_mul_componentxUMxa4_and_b9,
         input_p1_times_b1_mul_componentxUMxa3_and_b10,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831568_127845824_127847728,
         input_p1_times_b1_mul_componentxUMxa2_and_b11,
         input_p1_times_b1_mul_componentxUMxa1_and_b12,
         input_p1_times_b1_mul_componentxUMxa0_and_b13,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127635920_127637824_127713520,
         input_p1_times_b1_mul_componentxUMxa11_and_b1,
         input_p1_times_b1_mul_componentxUMxa10_and_b2,
         input_p1_times_b1_mul_componentxUMxa9_and_b3,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732480_127722160_127724064,
         input_p1_times_b1_mul_componentxUMxa8_and_b4,
         input_p1_times_b1_mul_componentxUMxa7_and_b5,
         input_p1_times_b1_mul_componentxUMxa6_and_b6,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673456_127675360_127730576,
         input_p1_times_b1_mul_componentxUMxa5_and_b7,
         input_p1_times_b1_mul_componentxUMxa4_and_b8,
         input_p1_times_b1_mul_componentxUMxa3_and_b9,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831456_127845712_127847616,
         input_p1_times_b1_mul_componentxUMxa2_and_b10,
         input_p1_times_b1_mul_componentxUMxa1_and_b11,
         input_p1_times_b1_mul_componentxUMxa0_and_b12,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127635808_127637712_127713408,
         input_p1_times_b1_mul_componentxUMxa11_and_b0,
         input_p1_times_b1_mul_componentxUMxa10_and_b1,
         input_p1_times_b1_mul_componentxUMxa9_and_b2,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732368_127722048_127723952,
         input_p1_times_b1_mul_componentxUMxa8_and_b3,
         input_p1_times_b1_mul_componentxUMxa7_and_b4,
         input_p1_times_b1_mul_componentxUMxa6_and_b5,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673344_127675248_127730464,
         input_p1_times_b1_mul_componentxUMxa5_and_b6,
         input_p1_times_b1_mul_componentxUMxa4_and_b7,
         input_p1_times_b1_mul_componentxUMxa3_and_b8,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831344_127845600_127847504,
         input_p1_times_b1_mul_componentxUMxa2_and_b9,
         input_p1_times_b1_mul_componentxUMxa1_and_b10,
         input_p1_times_b1_mul_componentxUMxa0_and_b11,
         input_p1_times_b1_mul_componentxUMxcarry_layer1_127635696_127637600,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127635696_127637600,
         input_p1_times_b1_mul_componentxUMxa10_and_b0,
         input_p1_times_b1_mul_componentxUMxa9_and_b1,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732256_127721936_127723840,
         input_p1_times_b1_mul_componentxUMxa8_and_b2,
         input_p1_times_b1_mul_componentxUMxa7_and_b3,
         input_p1_times_b1_mul_componentxUMxa6_and_b4,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673232_127675136_127730352,
         input_p1_times_b1_mul_componentxUMxa5_and_b5,
         input_p1_times_b1_mul_componentxUMxa4_and_b6,
         input_p1_times_b1_mul_componentxUMxa3_and_b7,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831232_127845488_127847392,
         input_p1_times_b1_mul_componentxUMxa2_and_b8,
         input_p1_times_b1_mul_componentxUMxa1_and_b9,
         input_p1_times_b1_mul_componentxUMxa0_and_b10,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732144_127721824_127723728,
         input_p1_times_b1_mul_componentxUMxa8_and_b1,
         input_p1_times_b1_mul_componentxUMxa7_and_b2,
         input_p1_times_b1_mul_componentxUMxa6_and_b3,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673120_127675024_127730240,
         input_p1_times_b1_mul_componentxUMxa5_and_b4,
         input_p1_times_b1_mul_componentxUMxa4_and_b5,
         input_p1_times_b1_mul_componentxUMxa3_and_b6,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831120_127845376_127847280,
         input_p1_times_b1_mul_componentxUMxa2_and_b7,
         input_p1_times_b1_mul_componentxUMxa1_and_b8,
         input_p1_times_b1_mul_componentxUMxa0_and_b9,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127732032_127721712_127723616,
         input_p1_times_b1_mul_componentxUMxa8_and_b0,
         input_p1_times_b1_mul_componentxUMxa7_and_b1,
         input_p1_times_b1_mul_componentxUMxa6_and_b2,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127673008_127674912_127730128,
         input_p1_times_b1_mul_componentxUMxa5_and_b3,
         input_p1_times_b1_mul_componentxUMxa4_and_b4,
         input_p1_times_b1_mul_componentxUMxa3_and_b5,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127831008_127845264_127847168,
         input_p1_times_b1_mul_componentxUMxa2_and_b6,
         input_p1_times_b1_mul_componentxUMxa1_and_b7,
         input_p1_times_b1_mul_componentxUMxa0_and_b8,
         input_p1_times_b1_mul_componentxUMxcarry_layer1_127731920_127721600,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127731920_127721600,
         input_p1_times_b1_mul_componentxUMxa7_and_b0,
         input_p1_times_b1_mul_componentxUMxa6_and_b1,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127672896_127674800_127730016,
         input_p1_times_b1_mul_componentxUMxa5_and_b2,
         input_p1_times_b1_mul_componentxUMxa4_and_b3,
         input_p1_times_b1_mul_componentxUMxa3_and_b4,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127830896_127845152_127847056,
         input_p1_times_b1_mul_componentxUMxa2_and_b5,
         input_p1_times_b1_mul_componentxUMxa1_and_b6,
         input_p1_times_b1_mul_componentxUMxa0_and_b7,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127672784_127674688_127729904,
         input_p1_times_b1_mul_componentxUMxa5_and_b1,
         input_p1_times_b1_mul_componentxUMxa4_and_b2,
         input_p1_times_b1_mul_componentxUMxa3_and_b3,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127830784_127845040_127846944,
         input_p1_times_b1_mul_componentxUMxa2_and_b4,
         input_p1_times_b1_mul_componentxUMxa1_and_b5,
         input_p1_times_b1_mul_componentxUMxa0_and_b6,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127672672_127674576_127729792,
         input_p1_times_b1_mul_componentxUMxa5_and_b0,
         input_p1_times_b1_mul_componentxUMxa4_and_b1,
         input_p1_times_b1_mul_componentxUMxa3_and_b2,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127830672_127844928_127846832,
         input_p1_times_b1_mul_componentxUMxa2_and_b3,
         input_p1_times_b1_mul_componentxUMxa1_and_b4,
         input_p1_times_b1_mul_componentxUMxa0_and_b5,
         input_p1_times_b1_mul_componentxUMxcarry_layer1_127672560_127674464,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127672560_127674464,
         input_p1_times_b1_mul_componentxUMxa4_and_b0,
         input_p1_times_b1_mul_componentxUMxa3_and_b1,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127830560_127844816_127846720,
         input_p1_times_b1_mul_componentxUMxa2_and_b2,
         input_p1_times_b1_mul_componentxUMxa1_and_b3,
         input_p1_times_b1_mul_componentxUMxa0_and_b4,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127830448_127844704_127846608,
         input_p1_times_b1_mul_componentxUMxa2_and_b1,
         input_p1_times_b1_mul_componentxUMxa1_and_b2,
         input_p1_times_b1_mul_componentxUMxa0_and_b3,
         input_p1_times_b1_mul_componentxUMxsum_layer1_127830336_127844592_127846496,
         input_p1_times_b1_mul_componentxUMxa2_and_b0,
         input_p1_times_b1_mul_componentxUMxa1_and_b1,
         input_p1_times_b1_mul_componentxUMxa0_and_b2,
         input_p1_times_b1_mul_componentxUMxcarry_layer1_127830168_127844480,
         input_p1_times_b1_mul_componentxUMxa1_and_b0,
         input_p1_times_b1_mul_componentxUMxa0_and_b1,
         output_p2_times_a2_div_componentxUDxis_less_than,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_0,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_1,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_2,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_3,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_4,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_5,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_6,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_7,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_8,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_9,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_10,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_11,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_12,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_13,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_14,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_15,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_16,
         output_p2_times_a2_div_componentxUDxcentral_parallel_output_17,
         output_p2_times_a2_div_componentxUDxshifted_substraction_result_0,
         output_p1_times_a1_div_componentxUDxis_less_than,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_0,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_1,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_2,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_3,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_4,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_5,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_6,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_7,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_8,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_9,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_10,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_11,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_12,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_13,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_14,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_15,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_16,
         output_p1_times_a1_div_componentxUDxcentral_parallel_output_17,
         output_p1_times_a1_div_componentxUDxshifted_substraction_result_0,
         input_p2_times_b2_div_componentxUDxis_less_than,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_0,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_1,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_2,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_3,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_4,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_5,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_6,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_7,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_8,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_9,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_10,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_11,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_12,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_13,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_14,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_15,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_16,
         input_p2_times_b2_div_componentxUDxcentral_parallel_output_17,
         input_p2_times_b2_div_componentxUDxshifted_substraction_result_0,
         input_p1_times_b1_div_componentxUDxis_less_than,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_0,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_1,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_2,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_3,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_4,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_5,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_6,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_7,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_8,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_9,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_10,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_11,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_12,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_13,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_14,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_15,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_16,
         input_p1_times_b1_div_componentxUDxcentral_parallel_output_17,
         input_p1_times_b1_div_componentxUDxshifted_substraction_result_0,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_0,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_1,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_2,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_3,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_4,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_5,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_6,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_7,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_8,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_9,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_10,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_11,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_12,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_13,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_14,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_15,
         output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_16,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_0,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_1,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_2,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_3,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_4,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_5,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_6,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_7,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_8,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_9,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_10,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_11,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_12,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_13,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_14,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_15,
         output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_16,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_0,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_1,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_2,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_3,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_4,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_5,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_6,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_7,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_8,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_9,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_10,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_11,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_12,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_13,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_14,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_15,
         input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_16,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_0,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_1,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_2,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_3,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_4,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_5,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_6,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_7,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_8,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_9,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_10,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_11,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_12,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_13,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_14,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_15,
         input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_16,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672;
  wire   [17:1] input_previous_0;
  wire   [17:1] input_previous_1;
  wire   [17:1] input_previous_2;
  wire   [17:8] output_previous_1;
  wire   [17:1] output_previous_2;
  wire   [17:0] results_b0_b1;
  wire   [17:0] results_b0_b1_b2;
  wire   [17:1] results_a1_a2;
  wire   [17:0] results_a1_a2_inv;
  wire   [17:1] input_times_b0_mul_componentxunsigned_output_inverted;
  wire   [17:0] input_times_b0_mul_componentxinput_A_inverted;
  wire   [17:0] input_times_b0_div_componentxunsigned_output_inverted;
  wire   [17:1] input_times_b0_div_componentxinput_A_inverted;
  wire   [21:0] clock_chopper_and_divisionxdivision_ring;
  wire   [17:7] input_times_b0_mul_componentxUMxsecond_vector;
  wire   [15:0] input_times_b0_mul_componentxUMxfirst_vector;
  wire   [18:0] input_times_b0_div_componentxUDxreadiness_propagation_vector;
  wire   [16:0] input_times_b0_div_componentxUDxsubstraction_result_too_long;
  wire   [16:1] input_times_b0_div_componentxUDxsub_ready_negative_divisor;
  wire   [17:0] input_times_b0_div_componentxUDxquotient_not_gated;
  wire   [17:1] output_p2_times_a2_mul_componentxunsigned_output_inverted;
  wire   [17:0] output_p2_times_a2_mul_componentxinput_A_inverted;
  wire   [17:1] output_p1_times_a1_mul_componentxunsigned_output_inverted;
  wire   [17:1] input_p2_times_b2_mul_componentxunsigned_output_inverted;
  wire   [17:0] input_p2_times_b2_mul_componentxinput_A_inverted;
  wire   [17:1] input_p1_times_b1_mul_componentxunsigned_output_inverted;
  wire   [17:0] input_p1_times_b1_mul_componentxinput_A_inverted;
  wire   [17:0] output_p2_times_a2_div_componentxunsigned_output_inverted;
  wire   [17:1] output_p2_times_a2_div_componentxinput_A_inverted;
  wire   [17:0] output_p1_times_a1_div_componentxunsigned_output_inverted;
  wire   [17:1] output_p1_times_a1_div_componentxinput_A_inverted;
  wire   [17:0] input_p2_times_b2_div_componentxunsigned_output_inverted;
  wire   [17:1] input_p2_times_b2_div_componentxinput_A_inverted;
  wire   [17:0] input_p1_times_b1_div_componentxunsigned_output_inverted;
  wire   [17:1] input_p1_times_b1_div_componentxinput_A_inverted;
  wire   [17:7] output_p2_times_a2_mul_componentxUMxsecond_vector;
  wire   [15:0] output_p2_times_a2_mul_componentxUMxfirst_vector;
  wire   [17:7] output_p1_times_a1_mul_componentxUMxsecond_vector;
  wire   [15:0] output_p1_times_a1_mul_componentxUMxfirst_vector;
  wire   [17:7] input_p2_times_b2_mul_componentxUMxsecond_vector;
  wire   [15:0] input_p2_times_b2_mul_componentxUMxfirst_vector;
  wire   [17:7] input_p1_times_b1_mul_componentxUMxsecond_vector;
  wire   [15:0] input_p1_times_b1_mul_componentxUMxfirst_vector;
  wire  
         [18:0] output_p2_times_a2_div_componentxUDxreadiness_propagation_vector
;
  wire  
         [16:0] output_p2_times_a2_div_componentxUDxsubstraction_result_too_long
;
  wire   [16:1] output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor
;
  wire   [17:0] output_p2_times_a2_div_componentxUDxquotient_not_gated;
  wire  
         [18:0] output_p1_times_a1_div_componentxUDxreadiness_propagation_vector
;
  wire  
         [16:0] output_p1_times_a1_div_componentxUDxsubstraction_result_too_long
;
  wire   [16:1] output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor
;
  wire   [17:0] output_p1_times_a1_div_componentxUDxquotient_not_gated;
  wire  
         [18:0] input_p2_times_b2_div_componentxUDxreadiness_propagation_vector
;
  wire  
         [16:0] input_p2_times_b2_div_componentxUDxsubstraction_result_too_long
;
  wire   [16:1] input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor;
  wire   [17:0] input_p2_times_b2_div_componentxUDxquotient_not_gated;
  wire  
         [18:0] input_p1_times_b1_div_componentxUDxreadiness_propagation_vector
;
  wire  
         [16:0] input_p1_times_b1_div_componentxUDxsubstraction_result_too_long
;
  wire   [16:1] input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor;
  wire   [17:0] input_p1_times_b1_div_componentxUDxquotient_not_gated;

  XOR2X4 final_adderxU53 ( .A(results_a1_a2_inv[0]), .B(results_b0_b1_b2[0]), 
        .Y(\output_signal[0] ) );
  XOR2X4 final_adderxU9 ( .A(n4166), .B(n4167), .Y(\output_signal[2] ) );
  XOR2X4 final_adderxU8 ( .A(n4164), .B(n4165), .Y(\output_signal[3] ) );
  XOR2X4 final_adderxU7 ( .A(n4162), .B(n4163), .Y(\output_signal[4] ) );
  XOR2X4 final_adderxU6 ( .A(n4160), .B(n4161), .Y(\output_signal[5] ) );
  XOR2X4 final_adderxU5 ( .A(n4158), .B(n4159), .Y(\output_signal[6] ) );
  XOR2X4 final_adderxU4 ( .A(n4156), .B(n4157), .Y(\output_signal[7] ) );
  DFFSX1 clock_chopper_and_divisionxdivision_ring_reg_1 ( 
        .D(clock_chopper_and_divisionxn47), .CK(clk), .SN(n283), 
        .Q(clock_chopper_and_divisionxdivision_ring[1]), .QN(n1261) );
  DFFSX1 clock_chopper_and_divisionxdivision_ring_reg_0 ( 
        .D(clock_chopper_and_divisionxn49), .CK(clk), .SN(n283), 
        .Q(clock_chopper_and_divisionxdivision_ring[0]), .QN(n1262) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_21 ( 
        .D(clock_chopper_and_divisionxn26), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[21]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_20 ( 
        .D(clock_chopper_and_divisionxn27), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[20]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_19 ( 
        .D(clock_chopper_and_divisionxn28), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[19]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_18 ( 
        .D(clock_chopper_and_divisionxn29), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[18]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_17 ( 
        .D(clock_chopper_and_divisionxn30), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[17]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_16 ( 
        .D(clock_chopper_and_divisionxn31), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[16]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_15 ( 
        .D(clock_chopper_and_divisionxn32), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[15]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_14 ( 
        .D(clock_chopper_and_divisionxn33), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[14]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_13 ( 
        .D(clock_chopper_and_divisionxn34), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[13]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_12 ( 
        .D(clock_chopper_and_divisionxn35), .CK(clk), .RN(n305), 
        .Q(clock_chopper_and_divisionxdivision_ring[12]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_11 ( 
        .D(clock_chopper_and_divisionxn36), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[11]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_10 ( 
        .D(clock_chopper_and_divisionxn37), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[10]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_9 ( 
        .D(clock_chopper_and_divisionxn38), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[9]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_8 ( 
        .D(clock_chopper_and_divisionxn39), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[8]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_7 ( 
        .D(clock_chopper_and_divisionxn40), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[7]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_6 ( 
        .D(clock_chopper_and_divisionxn41), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[6]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_5 ( 
        .D(clock_chopper_and_divisionxn42), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[5]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_4 ( 
        .D(clock_chopper_and_divisionxn43), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[4]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_3 ( 
        .D(clock_chopper_and_divisionxn44), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[3]) );
  DFFRHQX1 clock_chopper_and_divisionxdivision_ring_reg_2 ( 
        .D(clock_chopper_and_divisionxn45), .CK(clk), .RN(n304), 
        .Q(clock_chopper_and_divisionxdivision_ring[2]) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_16 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn23), .CK(clk), 
        .RN(n302), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_16) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_15 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn24), .CK(clk), 
        .RN(n302), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_15) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_14 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn25), .CK(clk), 
        .RN(n302), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_14) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_13 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn26), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_13) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_12 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn27), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_12) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_11 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn28), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_11) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_10 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn29), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_10) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_9 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn30), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_9) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_8 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn31), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_8) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_7 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn32), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_7) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_6 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn33), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_6) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_5 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn34), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_5) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_4 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn35), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_4) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_3 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn36), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_3) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_2 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn37), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_2) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_1 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn38), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_1) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_0 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn40), .CK(clk), 
        .RN(n301), 
        .Q(input_times_b0_div_componentxUDxinput_containerxparallel_out_0) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_16 ( 
        .D(n2218), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_16)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_15 ( 
        .D(n2219), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_15)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_14 ( 
        .D(n2220), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_14)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_13 ( 
        .D(n2221), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_13)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_12 ( 
        .D(n2222), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_12)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_11 ( 
        .D(n2223), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_11)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_10 ( 
        .D(n2224), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_10)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_9 ( 
        .D(n2225), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_9)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_8 ( 
        .D(n2226), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_8)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_7 ( 
        .D(n2227), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_7)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_6 ( 
        .D(n2228), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_6)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_5 ( 
        .D(n2229), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_5)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_4 ( 
        .D(n2230), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_4)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_3 ( 
        .D(n2231), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_3)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_2 ( 
        .D(n2232), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_2)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_1 ( 
        .D(n2233), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_1)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_0 ( 
        .D(n2234), .CK(clk), .RN(n286), 
        .Q(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_0)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_16 ( 
        .D(n2109), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_16)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_15 ( 
        .D(n2110), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_15)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_14 ( 
        .D(n2111), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_14)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_13 ( 
        .D(n2112), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_13)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_12 ( 
        .D(n2113), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_12)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_11 ( 
        .D(n2114), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_11)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_10 ( 
        .D(n2115), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_10)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_9 ( 
        .D(n2116), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_9)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_8 ( 
        .D(n2117), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_8)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_7 ( 
        .D(n2118), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_7)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_6 ( 
        .D(n2119), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_6)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_5 ( 
        .D(n2120), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_5)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_4 ( 
        .D(n2121), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_4)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_3 ( 
        .D(n2122), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_3)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_2 ( 
        .D(n2123), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_2)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_1 ( 
        .D(n2124), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_1)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_0 ( 
        .D(n2125), .CK(clk), .RN(n283), 
        .Q(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_0)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_16 ( 
        .D(n1999), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_16)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_15 ( 
        .D(n2000), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_15)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_14 ( 
        .D(n2001), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_14)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_13 ( 
        .D(n2002), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_13)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_12 ( 
        .D(n2003), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_12)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_11 ( 
        .D(n2004), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_11)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_10 ( 
        .D(n2005), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_10)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_9 ( 
        .D(n2006), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_9)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_8 ( 
        .D(n2007), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_8)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_7 ( 
        .D(n2008), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_7)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_6 ( 
        .D(n2009), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_6)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_5 ( 
        .D(n2010), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_5)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_4 ( 
        .D(n2011), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_4)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_3 ( 
        .D(n2012), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_3)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_2 ( 
        .D(n2013), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_2)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_1 ( 
        .D(n2014), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_1)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_0 ( 
        .D(n2015), .CK(clk), .RN(n295), 
        .Q(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_0)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_16 ( 
        .D(n1890), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_16)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_15 ( 
        .D(n1891), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_15)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_14 ( 
        .D(n1892), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_14)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_13 ( 
        .D(n1893), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_13)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_12 ( 
        .D(n1894), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_12)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_11 ( 
        .D(n1895), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_11)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_10 ( 
        .D(n1896), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_10)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_9 ( 
        .D(n1897), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_9)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_8 ( 
        .D(n1898), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_8)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_7 ( 
        .D(n1899), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_7)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_6 ( 
        .D(n1900), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_6)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_5 ( 
        .D(n1901), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_5)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_4 ( 
        .D(n1902), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_4)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_3 ( 
        .D(n1903), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_3)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_2 ( 
        .D(n1904), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_2)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_1 ( 
        .D(n1905), .CK(clk), .RN(n292), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_1)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_0 ( 
        .D(n1906), .CK(clk), .RN(n292), 
        .Q(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_0)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_19 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[18]), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxoutput_ready_signal) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_19 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[18]), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxoutput_ready_signal) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_19 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[18]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxoutput_ready_signal) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_17 ( 
        .D(n2289), .CK(clk), .RN(n289), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[17]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_17 ( 
        .D(n2180), .CK(clk), .RN(n286), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[17]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_17 ( 
        .D(n2070), .CK(clk), .RN(n283), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[17]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_17 ( 
        .D(n1961), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[17]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_17 ( 
        .D(n1851), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[17]) );
  DFFRHQX1 input_times_b0_div_componentxoutput_sign_gated_prev_reg ( .D(n379), 
        .CK(clk), .RN(n305), 
        .Q(input_times_b0_div_componentxoutput_sign_gated_prev) );
  DFFRHQX1 output_p2_times_a2_div_componentxoutput_sign_gated_prev_reg ( 
        .D(n377), .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxoutput_sign_gated_prev) );
  DFFRHQX1 input_p2_times_b2_div_componentxoutput_sign_gated_prev_reg ( 
        .D(n375), .CK(clk), .RN(n313), 
        .Q(input_p2_times_b2_div_componentxoutput_sign_gated_prev) );
  DFFRHQX1 input_p1_times_b1_div_componentxoutput_sign_gated_prev_reg ( 
        .D(n373), .CK(clk), .RN(n313), 
        .Q(input_p1_times_b1_div_componentxoutput_sign_gated_prev) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_16 ( 
        .D(n2290), .CK(clk), .RN(n289), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[16]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_15 ( 
        .D(n2291), .CK(clk), .RN(n289), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[15]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_14 ( 
        .D(n2292), .CK(clk), .RN(n289), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[14]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_13 ( 
        .D(n2293), .CK(clk), .RN(n289), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[13]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_12 ( 
        .D(n2294), .CK(clk), .RN(n289), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[12]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_11 ( 
        .D(n2295), .CK(clk), .RN(n289), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[11]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_10 ( 
        .D(n2296), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[10]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_9 ( 
        .D(n2297), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[9]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_8 ( 
        .D(n2298), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[8]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_7 ( 
        .D(n2299), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[7]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_6 ( 
        .D(n2300), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[6]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_5 ( 
        .D(n2301), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[5]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_4 ( 
        .D(n2302), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[4]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_3 ( 
        .D(n2303), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[3]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_2 ( 
        .D(n2304), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[2]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_1 ( 
        .D(n2305), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[1]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_0 ( 
        .D(n2306), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxquotient_not_gated[0]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_16 ( 
        .D(n2181), .CK(clk), .RN(n286), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[16]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_15 ( 
        .D(n2182), .CK(clk), .RN(n286), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[15]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_14 ( 
        .D(n2183), .CK(clk), .RN(n286), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[14]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_13 ( 
        .D(n2184), .CK(clk), .RN(n286), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[13]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_12 ( 
        .D(n2185), .CK(clk), .RN(n286), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[12]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_11 ( 
        .D(n2186), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[11]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_10 ( 
        .D(n2187), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[10]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_9 ( 
        .D(n2188), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[9]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_8 ( 
        .D(n2189), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[8]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_7 ( 
        .D(n2190), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[7]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_6 ( 
        .D(n2191), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[6]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_5 ( 
        .D(n2192), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[5]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_4 ( 
        .D(n2193), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[4]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_3 ( 
        .D(n2194), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[3]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_2 ( 
        .D(n2195), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[2]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_1 ( 
        .D(n2196), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[1]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_0 ( 
        .D(n2197), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxquotient_not_gated[0]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_16 ( 
        .D(n2071), .CK(clk), .RN(n283), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[16]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_15 ( 
        .D(n2072), .CK(clk), .RN(n287), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[15]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_14 ( 
        .D(n2073), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[14]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_13 ( 
        .D(n2074), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[13]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_12 ( 
        .D(n2075), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[12]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_11 ( 
        .D(n2076), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[11]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_10 ( 
        .D(n2077), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[10]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_9 ( 
        .D(n2078), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[9]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_8 ( 
        .D(n2079), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[8]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_7 ( 
        .D(n2080), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[7]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_6 ( 
        .D(n2081), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[6]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_5 ( 
        .D(n2082), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[5]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_4 ( 
        .D(n2083), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[4]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_3 ( 
        .D(n2084), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[3]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_2 ( 
        .D(n2085), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[2]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_1 ( 
        .D(n2086), .CK(clk), .RN(n298), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[1]) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_0 ( 
        .D(n2087), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxquotient_not_gated[0]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_16 ( 
        .D(n1962), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[16]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_15 ( 
        .D(n1963), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[15]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_14 ( 
        .D(n1964), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[14]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_13 ( 
        .D(n1965), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[13]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_12 ( 
        .D(n1966), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[12]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_11 ( 
        .D(n1967), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[11]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_10 ( 
        .D(n1968), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[10]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_9 ( 
        .D(n1969), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[9]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_8 ( 
        .D(n1970), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[8]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_7 ( 
        .D(n1971), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[7]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_6 ( 
        .D(n1972), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[6]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_5 ( 
        .D(n1973), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[5]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_4 ( 
        .D(n1974), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[4]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_3 ( 
        .D(n1975), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[3]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_2 ( 
        .D(n1976), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[2]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_1 ( 
        .D(n1977), .CK(clk), .RN(n295), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[1]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_0 ( 
        .D(n1978), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxquotient_not_gated[0]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_16 ( 
        .D(n1852), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[16]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_15 ( 
        .D(n1853), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[15]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_14 ( 
        .D(n1854), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[14]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_13 ( 
        .D(n1855), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[13]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_12 ( 
        .D(n1856), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[12]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_11 ( 
        .D(n1857), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[11]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_10 ( 
        .D(n1858), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[10]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_9 ( 
        .D(n1859), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[9]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_8 ( 
        .D(n1860), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[8]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_7 ( 
        .D(n1861), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[7]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_6 ( 
        .D(n1862), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[6]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_5 ( 
        .D(n1863), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[5]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_4 ( 
        .D(n1864), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[4]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_3 ( 
        .D(n1865), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[3]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_2 ( 
        .D(n1866), .CK(clk), .RN(n292), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[2]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_1 ( 
        .D(n1867), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[1]) );
  DFFRHQX1 input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_0 ( 
        .D(n1868), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxquotient_not_gated[0]) );
  DFFRHQX1 input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_17 ( 
        .D(input_times_b0_div_componentxUDxinput_containerxn22), .CK(clk), 
        .RN(n302), 
        .Q(input_times_b0_div_componentxUDxshifted_substraction_result_0) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_17 ( 
        .D(n2217), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxshifted_substraction_result_0)
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_17 ( 
        .D(n2108), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxshifted_substraction_result_0)
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_17 ( 
        .D(n1998), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxshifted_substraction_result_0)
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_17 ( 
        .D(n1889), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxshifted_substraction_result_0)
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_17 ( 
        .D(n2253), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_17) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_17 ( 
        .D(n2144), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_17) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_17 ( 
        .D(n2034), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_17) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_17 ( 
        .D(n1925), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_17) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_17 ( 
        .D(n1815), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_17) );
  DFFRHQX1 clock_chopper_and_divisionxclk_out_reg ( 
        .D(clock_chopper_and_divisionxn46), .CK(clk), .RN(n304), .Q(n4673) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_16 ( 
        .D(n2254), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_16) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_16 ( 
        .D(n2145), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_16) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_16 ( 
        .D(n2035), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_16) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_16 ( 
        .D(n1926), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_16) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_16 ( 
        .D(n1816), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_16) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_14 ( 
        .D(n2256), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_14) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_14 ( 
        .D(n2147), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_14) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_14 ( 
        .D(n2037), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_14) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_14 ( 
        .D(n1928), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_14) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_14 ( 
        .D(n1818), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_14) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_15 ( 
        .D(n2255), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_15) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_15 ( 
        .D(n2146), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_15) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_15 ( 
        .D(n2036), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_15) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_15 ( 
        .D(n1927), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_15) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_15 ( 
        .D(n1817), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_15) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_12 ( 
        .D(n2258), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_12) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_10 ( 
        .D(n2260), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_10) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_8 ( 
        .D(n2262), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_8) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_12 ( 
        .D(n2149), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_12) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_10 ( 
        .D(n2151), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_10) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_8 ( 
        .D(n2153), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_8) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_12 ( 
        .D(n2039), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_12) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_10 ( 
        .D(n2041), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_10) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_8 ( 
        .D(n2043), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_8) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_12 ( 
        .D(n1930), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_12) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_10 ( 
        .D(n1932), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_10) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_8 ( 
        .D(n1934), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_8) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_12 ( 
        .D(n1820), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_12) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_10 ( 
        .D(n1822), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_10) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_8 ( 
        .D(n1824), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_8) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_13 ( 
        .D(n2257), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_13) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_11 ( 
        .D(n2259), .CK(clk), .RN(n288), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_11) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_9 ( 
        .D(n2261), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_9) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_13 ( 
        .D(n2148), .CK(clk), .RN(n285), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_13) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_11 ( 
        .D(n2150), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_11) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_9 ( 
        .D(n2152), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_9) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_13 ( 
        .D(n2038), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_13) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_11 ( 
        .D(n2040), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_11) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_9 ( 
        .D(n2042), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_9) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_13 ( 
        .D(n1929), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_13) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_11 ( 
        .D(n1931), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_11) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_9 ( 
        .D(n1933), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_9) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_13 ( 
        .D(n1819), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_13) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_11 ( 
        .D(n1821), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_11) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_9 ( 
        .D(n1823), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_9) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_6 ( 
        .D(n2264), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_6) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_4 ( 
        .D(n2266), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_4) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_6 ( 
        .D(n2155), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_6) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_4 ( 
        .D(n2157), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_4) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_6 ( 
        .D(n2045), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_6) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_4 ( 
        .D(n2047), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_4) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_6 ( 
        .D(n1936), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_6) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_4 ( 
        .D(n1938), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_4) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_6 ( 
        .D(n1826), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_6) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_4 ( 
        .D(n1828), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_4) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_7 ( 
        .D(n2263), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_7) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_5 ( 
        .D(n2265), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_5) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_7 ( 
        .D(n2154), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_7) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_5 ( 
        .D(n2156), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_5) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_7 ( 
        .D(n2044), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_7) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_5 ( 
        .D(n2046), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_5) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_7 ( 
        .D(n1935), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_7) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_5 ( 
        .D(n1937), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_5) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_7 ( 
        .D(n1825), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_7) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_5 ( 
        .D(n1827), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_5) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_2 ( 
        .D(n2268), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_2) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_2 ( 
        .D(n2159), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_2) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_2 ( 
        .D(n2049), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_2) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_2 ( 
        .D(n1940), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_2) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_2 ( 
        .D(n1830), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_2) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_0 ( 
        .D(n2270), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_0) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_0 ( 
        .D(n2161), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_0) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_0 ( 
        .D(n2051), .CK(clk), .RN(n296), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_0) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_0 ( 
        .D(n1942), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_0) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_0 ( 
        .D(n1832), .CK(clk), .RN(n298), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_0) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_1 ( 
        .D(n2269), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_1) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_1 ( 
        .D(n2160), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_1) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_1 ( 
        .D(n2050), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_1) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_1 ( 
        .D(n1941), .CK(clk), .RN(n293), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_1) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_1 ( 
        .D(n1831), .CK(clk), .RN(n294), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_1) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_3 ( 
        .D(n2267), .CK(clk), .RN(n287), 
        .Q(output_p2_times_a2_div_componentxUDxcentral_parallel_output_3) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_3 ( 
        .D(n2158), .CK(clk), .RN(n284), 
        .Q(output_p1_times_a1_div_componentxUDxcentral_parallel_output_3) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_3 ( 
        .D(n2048), .CK(clk), .RN(n297), 
        .Q(input_p2_times_b2_div_componentxUDxcentral_parallel_output_3) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_3 ( 
        .D(n1939), .CK(clk), .RN(n294), 
        .Q(input_p1_times_b1_div_componentxUDxcentral_parallel_output_3) );
  DFFRHQX1 input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_3 ( 
        .D(n1829), .CK(clk), .RN(n291), 
        .Q(input_times_b0_div_componentxUDxcentral_parallel_output_3) );
  DFFRHQX1 output_prev_2_registerxq_reg_16 ( .D(n4671), .CK(clk), .RN(n300), 
        .Q(output_previous_2[16]) );
  DFFRHQX1 input_prev_2_registerxq_reg_16 ( .D(n4653), .CK(clk), .RN(n299), 
        .Q(input_previous_2[16]) );
  DFFRHQX1 output_prev_2_registerxq_reg_14 ( .D(n4669), .CK(clk), .RN(n300), 
        .Q(output_previous_2[14]) );
  DFFRHQX1 input_prev_2_registerxq_reg_14 ( .D(n4651), .CK(clk), .RN(n299), 
        .Q(input_previous_2[14]) );
  DFFRHQX1 output_prev_2_registerxq_reg_15 ( .D(n4670), .CK(clk), .RN(n300), 
        .Q(output_previous_2[15]) );
  DFFRHQX1 input_prev_2_registerxq_reg_15 ( .D(n4652), .CK(clk), .RN(n299), 
        .Q(input_previous_2[15]) );
  DFFRHQX1 input_prev_0_registerxq_reg_16 ( .D(input_prev_0_registerxn18), 
        .CK(clk), .RN(n305), .Q(input_previous_0[16]) );
  DFFRHQX1 input_prev_1_registerxq_reg_16 ( .D(n4635), .CK(clk), .RN(n313), 
        .Q(input_previous_1[16]) );
  DFFRHQX1 input_prev_0_registerxq_reg_15 ( .D(input_prev_0_registerxn17), 
        .CK(clk), .RN(n305), .Q(input_previous_0[15]) );
  DFFRHQX1 input_prev_1_registerxq_reg_15 ( .D(n4634), .CK(clk), .RN(n313), 
        .Q(input_previous_1[15]) );
  DFFRHQX1 output_prev_2_registerxq_reg_12 ( .D(n4667), .CK(clk), .RN(n300), 
        .Q(output_previous_2[12]) );
  DFFRHQX1 input_prev_2_registerxq_reg_12 ( .D(n4649), .CK(clk), .RN(n299), 
        .Q(input_previous_2[12]) );
  DFFRHQX1 output_prev_2_registerxq_reg_13 ( .D(n4668), .CK(clk), .RN(n300), 
        .Q(output_previous_2[13]) );
  DFFRHQX1 input_prev_2_registerxq_reg_13 ( .D(n4650), .CK(clk), .RN(n299), 
        .Q(input_previous_2[13]) );
  DFFRHQX1 input_prev_0_registerxq_reg_14 ( .D(input_prev_0_registerxn16), 
        .CK(clk), .RN(n305), .Q(input_previous_0[14]) );
  DFFRHQX1 input_prev_1_registerxq_reg_14 ( .D(n4633), .CK(clk), .RN(n314), 
        .Q(input_previous_1[14]) );
  DFFRHQX1 input_prev_0_registerxq_reg_13 ( .D(input_prev_0_registerxn15), 
        .CK(clk), .RN(n305), .Q(input_previous_0[13]) );
  DFFRHQX1 input_prev_1_registerxq_reg_13 ( .D(n4632), .CK(clk), .RN(n314), 
        .Q(input_previous_1[13]) );
  DFFRHQX1 output_prev_2_registerxq_reg_10 ( .D(n4665), .CK(clk), .RN(n300), 
        .Q(output_previous_2[10]) );
  DFFRHQX1 input_prev_2_registerxq_reg_10 ( .D(n4647), .CK(clk), .RN(n299), 
        .Q(input_previous_2[10]) );
  DFFRHQX1 output_prev_2_registerxq_reg_11 ( .D(n4666), .CK(clk), .RN(n300), 
        .Q(output_previous_2[11]) );
  DFFRHQX1 input_prev_2_registerxq_reg_11 ( .D(n4648), .CK(clk), .RN(n299), 
        .Q(input_previous_2[11]) );
  DFFRHQX1 input_prev_0_registerxq_reg_9 ( .D(input_prev_0_registerxn11), 
        .CK(clk), .RN(n306), .Q(input_previous_0[9]) );
  DFFRHQX1 output_prev_2_registerxq_reg_9 ( .D(n4664), .CK(clk), .RN(n300), 
        .Q(output_previous_2[9]) );
  DFFRHQX1 input_prev_2_registerxq_reg_9 ( .D(n4646), .CK(clk), .RN(n299), 
        .Q(input_previous_2[9]) );
  DFFRHQX1 input_prev_1_registerxq_reg_9 ( .D(n4628), .CK(clk), .RN(n314), 
        .Q(input_previous_1[9]) );
  DFFRHQX1 input_prev_0_registerxq_reg_10 ( .D(input_prev_0_registerxn12), 
        .CK(clk), .RN(n306), .Q(input_previous_0[10]) );
  DFFRHQX1 input_prev_1_registerxq_reg_10 ( .D(n4629), .CK(clk), .RN(n314), 
        .Q(input_previous_1[10]) );
  DFFRHQX1 input_prev_0_registerxq_reg_12 ( .D(input_prev_0_registerxn14), 
        .CK(clk), .RN(n305), .Q(input_previous_0[12]) );
  DFFRHQX1 input_prev_1_registerxq_reg_12 ( .D(n4631), .CK(clk), .RN(n314), 
        .Q(input_previous_1[12]) );
  DFFRHQX1 input_prev_0_registerxq_reg_11 ( .D(input_prev_0_registerxn13), 
        .CK(clk), .RN(n306), .Q(input_previous_0[11]) );
  DFFRHQX1 input_prev_1_registerxq_reg_11 ( .D(n4630), .CK(clk), .RN(n314), 
        .Q(input_previous_1[11]) );
  DFFRHQX1 input_prev_0_registerxq_reg_17 ( .D(input_prev_0_registerxn20), 
        .CK(clk), .RN(n305), .Q(input_previous_0[17]) );
  DFFRHQX1 output_prev_2_registerxq_reg_17 ( .D(n4672), .CK(clk), .RN(n300), 
        .Q(output_previous_2[17]) );
  DFFRHQX1 input_prev_2_registerxq_reg_17 ( .D(n4654), .CK(clk), .RN(n299), 
        .Q(input_previous_2[17]) );
  DFFRHQX1 input_prev_1_registerxq_reg_17 ( .D(n4636), .CK(clk), .RN(n313), 
        .Q(input_previous_1[17]) );
  DFFRHQX1 output_prev_2_registerxq_reg_4 ( .D(n4659), .CK(clk), .RN(n300), 
        .Q(output_previous_2[4]) );
  DFFRHQX1 output_prev_2_registerxq_reg_6 ( .D(n4661), .CK(clk), .RN(n300), 
        .Q(output_previous_2[6]) );
  DFFRHQX1 input_prev_2_registerxq_reg_4 ( .D(n4641), .CK(clk), .RN(n299), 
        .Q(input_previous_2[4]) );
  DFFRHQX1 input_prev_2_registerxq_reg_6 ( .D(n4643), .CK(clk), .RN(n299), 
        .Q(input_previous_2[6]) );
  DFFRHQX1 output_prev_2_registerxq_reg_8 ( .D(n4663), .CK(clk), .RN(n300), 
        .Q(output_previous_2[8]) );
  DFFRHQX1 input_prev_2_registerxq_reg_8 ( .D(n4645), .CK(clk), .RN(n299), 
        .Q(input_previous_2[8]) );
  DFFRHQX1 output_prev_2_registerxq_reg_3 ( .D(n4658), .CK(clk), .RN(n301), 
        .Q(output_previous_2[3]) );
  DFFRHQX1 output_prev_2_registerxq_reg_5 ( .D(n4660), .CK(clk), .RN(n300), 
        .Q(output_previous_2[5]) );
  DFFRHQX1 input_prev_2_registerxq_reg_3 ( .D(n4640), .CK(clk), .RN(n300), 
        .Q(input_previous_2[3]) );
  DFFRHQX1 input_prev_2_registerxq_reg_5 ( .D(n4642), .CK(clk), .RN(n299), 
        .Q(input_previous_2[5]) );
  DFFRHQX1 output_prev_2_registerxq_reg_7 ( .D(n4662), .CK(clk), .RN(n300), 
        .Q(output_previous_2[7]) );
  DFFRHQX1 input_prev_2_registerxq_reg_7 ( .D(n4644), .CK(clk), .RN(n299), 
        .Q(input_previous_2[7]) );
  DFFRHQX1 input_prev_0_registerxq_reg_4 ( .D(input_prev_0_registerxn6), 
        .CK(clk), .RN(n306), .Q(input_previous_0[4]) );
  DFFRHQX1 input_prev_0_registerxq_reg_6 ( .D(input_prev_0_registerxn8), 
        .CK(clk), .RN(n306), .Q(input_previous_0[6]) );
  DFFRHQX1 input_prev_1_registerxq_reg_4 ( .D(n4623), .CK(clk), .RN(n298), 
        .Q(input_previous_1[4]) );
  DFFRHQX1 input_prev_1_registerxq_reg_6 ( .D(n4625), .CK(clk), .RN(n298), 
        .Q(input_previous_1[6]) );
  DFFRHQX1 input_prev_0_registerxq_reg_8 ( .D(input_prev_0_registerxn10), 
        .CK(clk), .RN(n306), .Q(input_previous_0[8]) );
  DFFRHQX1 input_prev_1_registerxq_reg_8 ( .D(n4627), .CK(clk), .RN(n314), 
        .Q(input_previous_1[8]) );
  DFFRHQX1 input_prev_0_registerxq_reg_3 ( .D(input_prev_0_registerxn5), 
        .CK(clk), .RN(n306), .Q(input_previous_0[3]) );
  DFFRHQX1 input_prev_0_registerxq_reg_5 ( .D(input_prev_0_registerxn7), 
        .CK(clk), .RN(n306), .Q(input_previous_0[5]) );
  DFFRHQX1 input_prev_1_registerxq_reg_3 ( .D(n4622), .CK(clk), .RN(n299), 
        .Q(input_previous_1[3]) );
  DFFRHQX1 input_prev_1_registerxq_reg_5 ( .D(n4624), .CK(clk), .RN(n298), 
        .Q(input_previous_1[5]) );
  DFFRHQX1 input_prev_0_registerxq_reg_7 ( .D(input_prev_0_registerxn9), 
        .CK(clk), .RN(n306), .Q(input_previous_0[7]) );
  DFFRHQX1 input_prev_1_registerxq_reg_7 ( .D(n4626), .CK(clk), .RN(n302), 
        .Q(input_previous_1[7]) );
  DFFRHQX1 output_prev_2_registerxq_reg_2 ( .D(n4657), .CK(clk), .RN(n301), 
        .Q(output_previous_2[2]) );
  DFFRHQX1 input_prev_2_registerxq_reg_2 ( .D(n4639), .CK(clk), .RN(n300), 
        .Q(input_previous_2[2]) );
  DFFRHQX1 output_prev_2_registerxq_reg_1 ( .D(n4656), .CK(clk), .RN(n301), 
        .Q(output_previous_2[1]) );
  DFFRHQX1 input_prev_2_registerxq_reg_1 ( .D(n4638), .CK(clk), .RN(n300), 
        .Q(input_previous_2[1]) );
  DFFRHQX1 input_prev_0_registerxq_reg_2 ( .D(input_prev_0_registerxn4), 
        .CK(clk), .RN(n306), .Q(input_previous_0[2]) );
  DFFRHQX1 input_prev_1_registerxq_reg_2 ( .D(n4621), .CK(clk), .RN(n299), 
        .Q(input_previous_1[2]) );
  DFFRHQX1 input_prev_0_registerxq_reg_1 ( .D(input_prev_0_registerxn3), 
        .CK(clk), .RN(n306), .Q(input_previous_0[1]) );
  DFFRHQX1 input_prev_1_registerxq_reg_1 ( .D(n4620), .CK(clk), .RN(n299), 
        .Q(input_previous_1[1]) );
  DFFRHQX1 output_prev_2_registerxq_reg_0 ( .D(n4655), .CK(clk), .RN(n301), 
        .Q(output_p2_times_a2_mul_componentxinput_A_inverted[0]) );
  DFFRHQX1 input_prev_2_registerxq_reg_0 ( .D(n4637), .CK(clk), .RN(n300), 
        .Q(input_p2_times_b2_mul_componentxinput_A_inverted[0]) );
  DFFRHQX1 input_prev_0_registerxq_reg_0 ( .D(input_prev_0_registerxn2), 
        .CK(clk), .RN(n283), 
        .Q(input_times_b0_mul_componentxinput_A_inverted[0]) );
  DFFRHQX1 input_prev_1_registerxq_reg_0 ( .D(n4619), .CK(clk), .RN(n299), 
        .Q(input_p1_times_b1_mul_componentxinput_A_inverted[0]) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_17 ( .D(n1281), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_17) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_17 ( .D(n1400), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_17) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_17 ( .D(n1419), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_17) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_17 ( .D(n1438), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_17) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_17 ( .D(n1457), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_17) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_16 ( .D(n1399), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_16) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_16 ( .D(n1418), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_16) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_16 ( .D(n1437), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_16) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_16 ( .D(n1280), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_16) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_16 ( .D(n1456), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_16) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_12 ( .D(n1433), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_12) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_14 ( .D(n1278), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_14) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_14 ( .D(n1397), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_14) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_14 ( .D(n1416), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_14) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_14 ( .D(n1435), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_14) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_14 ( .D(n1454), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_14) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_15 ( .D(n1279), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_15) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_15 ( .D(n1398), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_15) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_15 ( .D(n1417), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_15) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_15 ( .D(n1436), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_15) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_15 ( .D(n1455), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_15) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_11 ( .D(n1432), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_11) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_13 ( .D(n1415), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_13) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_13 ( .D(n1434), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_13) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_10 ( .D(n1274), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_10) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_10 ( .D(n1393), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_10) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_10 ( .D(n1412), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_10) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_10 ( .D(n1431), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_10) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_10 ( .D(n1450), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_10) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_12 ( .D(n1276), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_12) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_12 ( .D(n1395), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_12) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_12 ( .D(n1414), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_12) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_12 ( .D(n1452), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_12) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_8 ( .D(n1428), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_8) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_11 ( .D(n1275), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_11) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_11 ( .D(n1394), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_11) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_11 ( .D(n1413), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_11) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_11 ( .D(n1451), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_11) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_9 ( .D(n1273), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_9) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_9 ( .D(n1392), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_9) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_9 ( .D(n1411), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_9) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_9 ( .D(n1430), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_9) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_13 ( .D(n1277), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_13) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_13 ( .D(n1396), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_13) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_7 ( .D(n1427), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_7) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_13 ( .D(n1453), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_13) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_2 ( .D(n1422), 
        .CK(clk), .RN(n309), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_2) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_6 ( .D(n1269), 
        .CK(clk), .RN(n304), 
        .Q(input_times_b0_div_componentxunsigned_output_6) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_6 ( .D(n1388), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_6) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_6 ( .D(n1407), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_6) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_4 ( .D(n1424), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_4) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_6 ( .D(n1426), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_6) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_6 ( .D(n1445), 
        .CK(clk), .RN(n306), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_6) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_8 ( .D(n1271), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_8) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_8 ( .D(n1390), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_8) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_8 ( .D(n1409), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_8) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_8 ( .D(n1447), 
        .CK(clk), .RN(n310), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_8) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_5 ( .D(n1268), 
        .CK(clk), .RN(n304), 
        .Q(input_times_b0_div_componentxunsigned_output_5) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_5 ( .D(n1387), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_5) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_5 ( .D(n1406), 
        .CK(clk), .RN(n311), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_5) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_3 ( .D(n1423), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_3) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_5 ( .D(n1425), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_5) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_5 ( .D(n1444), 
        .CK(clk), .RN(n306), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_5) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_9 ( .D(n1449), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_9) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_7 ( .D(n1270), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxunsigned_output_7) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_7 ( .D(n1389), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_7) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_7 ( .D(n1408), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_7) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_7 ( .D(n1446), 
        .CK(clk), .RN(n306), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_7) );
  DFFRHQX1 input_p2_times_b2_div_componentxoutput_sign_gated_reg ( .D(n4296), 
        .CK(clk), .RN(n313), 
        .Q(input_p2_times_b2_div_componentxoutput_sign_gated) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_2 ( .D(n1265), 
        .CK(clk), .RN(n304), 
        .Q(input_times_b0_div_componentxunsigned_output_2) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_2 ( .D(n1384), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_2) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_2 ( .D(n1403), 
        .CK(clk), .RN(n311), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_2) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_2 ( .D(n1441), 
        .CK(clk), .RN(n306), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_2) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_4 ( .D(n1267), 
        .CK(clk), .RN(n304), 
        .Q(input_times_b0_div_componentxunsigned_output_4) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_4 ( .D(n1386), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_4) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_4 ( .D(n1405), 
        .CK(clk), .RN(n311), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_4) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_4 ( .D(n1443), 
        .CK(clk), .RN(n306), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_4) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_1 ( .D(n1264), 
        .CK(clk), .RN(n304), 
        .Q(input_times_b0_div_componentxunsigned_output_1) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_1 ( .D(n1383), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_1) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_1 ( .D(n1402), 
        .CK(clk), .RN(n311), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_1) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_1 ( .D(n1421), 
        .CK(clk), .RN(n309), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_1) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_3 ( .D(n1266), 
        .CK(clk), .RN(n304), 
        .Q(input_times_b0_div_componentxunsigned_output_3) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_3 ( .D(n1385), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_3) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_3 ( .D(n1404), 
        .CK(clk), .RN(n311), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_3) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_3 ( .D(n1442), 
        .CK(clk), .RN(n306), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_3) );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxquotient_reg_0 ( .D(n1420), 
        .CK(clk), .RN(n309), 
        .Q(input_p2_times_b2_div_componentxunsigned_output_inverted[0]) );
  DFFRHQX1 input_times_b0_div_componentxoutput_sign_gated_reg ( 
        .D(input_times_b0_div_componentxn62), .CK(clk), .RN(n305), 
        .Q(input_times_b0_div_componentxoutput_sign_gated) );
  DFFRHQX1 output_p2_times_a2_div_componentxoutput_sign_gated_reg ( .D(n4406), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxoutput_sign_gated) );
  DFFRHQX1 output_p1_times_a1_div_componentxoutput_sign_gated_reg ( .D(n4350), 
        .CK(clk), .RN(n313), 
        .Q(output_p1_times_a1_div_componentxoutput_sign_gated) );
  DFFRHQX1 input_p1_times_b1_div_componentxoutput_sign_gated_reg ( .D(n4240), 
        .CK(clk), .RN(n313), 
        .Q(input_p1_times_b1_div_componentxoutput_sign_gated) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_1 ( .D(n1440), 
        .CK(clk), .RN(n306), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_1) );
  DFFRHQX1 input_times_b0_div_componentxUDxquotient_reg_0 ( .D(n1263), 
        .CK(clk), .RN(n304), 
        .Q(input_times_b0_div_componentxunsigned_output_inverted[0]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxquotient_reg_0 ( .D(n1382), 
        .CK(clk), .RN(n313), 
        .Q(output_p2_times_a2_div_componentxunsigned_output_inverted[0]) );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxquotient_reg_0 ( .D(n1401), 
        .CK(clk), .RN(n311), 
        .Q(output_p1_times_a1_div_componentxunsigned_output_inverted[0]) );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxquotient_reg_0 ( .D(n1439), 
        .CK(clk), .RN(n307), 
        .Q(input_p1_times_b1_div_componentxunsigned_output_inverted[0]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_0 ( 
        .D(change_input), .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[0]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_0 ( 
        .D(change_input), .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[0])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_0 ( 
        .D(change_input), .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[0])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_0 ( 
        .D(change_input), .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[0])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_0 ( 
        .D(change_input), .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[0])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_18 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[17]), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[18])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_17 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[16]), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[17])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_16 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[15]), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[16])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_15 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[14]), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[15])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_14 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[13]), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[14])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_13 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[12]), 
        .CK(clk), .RN(n303), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[13])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_12 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[11]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[12])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_11 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[10]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[11])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_10 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[9]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[10])
         );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_9 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[8]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[9]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_8 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[7]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[8]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_7 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[6]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[7]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_6 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[5]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[6]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_5 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[4]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[5]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_4 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[3]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[4]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_3 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[2]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[3]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_2 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[1]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[2]) );
  DFFRHQX1 input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_1 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[0]), 
        .CK(clk), .RN(n302), 
        .Q(input_times_b0_div_componentxUDxreadiness_propagation_vector[1]) );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_18 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[17]), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[18])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_17 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[16]), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[17])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_16 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[15]), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[16])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_15 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[14]), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[15])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_14 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[13]), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[14])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_13 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[12]), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[13])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_12 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[11]), 
        .CK(clk), .RN(n312), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[12])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_11 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[10]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[11])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_10 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[9]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[10])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_9 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[8]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[9])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_8 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[7]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[8])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_7 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[6]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[7])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_6 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[5]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[6])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_5 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[4]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[5])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_4 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[3]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[4])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_3 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[2]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[3])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_2 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[1]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[2])
         );
  DFFRHQX1 output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_1 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[0]), 
        .CK(clk), .RN(n311), 
        .Q(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[1])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_18 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[17]), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[18])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_17 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[16]), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[17])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_16 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[15]), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[16])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_15 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[14]), 
        .CK(clk), .RN(n310), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[15])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_14 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[13]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[14])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_13 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[12]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[13])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_12 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[11]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[12])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_11 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[10]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[11])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_10 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[9]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[10])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_9 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[8]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[9])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_8 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[7]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[8])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_7 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[6]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[7])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_6 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[5]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[6])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_5 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[4]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[5])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_4 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[3]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[4])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_3 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[2]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[3])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_2 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[1]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[2])
         );
  DFFRHQX1 output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_1 ( 
        .D(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[0]), 
        .CK(clk), .RN(n309), 
        .Q(output_p1_times_a1_div_componentxUDxreadiness_propagation_vector[1])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_18 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[17]), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[18])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_17 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[16]), 
        .CK(clk), .RN(n308), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[17])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_16 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[15]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[16])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_15 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[14]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[15])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_14 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[13]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[14])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_13 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[12]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[13])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_12 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[11]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[12])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_11 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[10]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[11])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_10 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[9]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[10])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_9 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[8]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[9])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_8 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[7]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[8])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_7 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[6]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[7])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_6 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[5]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[6])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_5 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[4]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[5])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_4 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[3]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[4])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_3 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[2]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[3])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_2 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[1]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[2])
         );
  DFFRHQX1 input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_1 ( 
        .D(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[0]), 
        .CK(clk), .RN(n307), 
        .Q(input_p2_times_b2_div_componentxUDxreadiness_propagation_vector[1])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_18 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[17]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[18])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_17 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[16]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[17])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_16 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[15]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[16])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_15 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[14]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[15])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_14 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[13]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[14])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_13 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[12]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[13])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_12 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[11]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[12])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_11 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[10]), 
        .CK(clk), .RN(n290), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[11])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_10 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[9]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[10])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_9 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[8]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[9])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_8 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[7]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[8])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_7 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[6]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[7])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_6 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[5]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[6])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_5 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[4]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[5])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_4 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[3]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[4])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_3 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[2]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[3])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_2 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[1]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[2])
         );
  DFFRHQX1 input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_1 ( 
        .D(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[0]), 
        .CK(clk), .RN(n289), 
        .Q(input_p1_times_b1_div_componentxUDxreadiness_propagation_vector[1])
         );
  DFFRXL input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_19 ( 
        .D(input_times_b0_div_componentxUDxreadiness_propagation_vector[18]), 
        .CK(clk), .RN(n283), .Q(n8), .QN(n257) );
  DFFRXL output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_19 ( 
        .D(output_p2_times_a2_div_componentxUDxreadiness_propagation_vector[18]), 
        .CK(clk), .RN(n284), .Q(n7), .QN(n164) );
  AND2X2 U3 ( .A(change_input), .B(en), .Y(n1) );
  NOR2X1 U4 ( .A(n367), .B(n837), .Y(n2) );
  NOR2X1 U5 ( .A(n368), .B(n996), .Y(n3) );
  NOR2X1 U6 ( .A(n367), .B(n1155), .Y(n4) );
  NOR2X1 U7 ( .A(n368), .B(n519), .Y(n5) );
  NOR2X1 U8 ( .A(n367), .B(n678), .Y(n6) );
  NAND2X1 U9 ( .A(output_p1_times_a1_mul_componentxinput_A_inverted_17_), 
        .B(n165), .Y(n9) );
  NAND2X1 U10 ( .A(input_p1_times_b1_mul_componentxinput_A_inverted[17]), 
        .B(input_previous_1[17]), .Y(n10) );
  NAND2X1 U11 ( .A(input_p2_times_b2_mul_componentxinput_A_inverted[17]), 
        .B(input_previous_2[17]), .Y(n11) );
  NAND2X1 U12 ( .A(output_p2_times_a2_mul_componentxinput_A_inverted[17]), 
        .B(output_previous_2[17]), .Y(n12) );
  NAND2X1 U13 ( .A(input_times_b0_mul_componentxinput_A_inverted[17]), 
        .B(input_previous_0[17]), .Y(n13) );
  AND2X2 U14 ( .A(n837), .B(en), .Y(n14) );
  AND2X2 U15 ( .A(n996), .B(en), .Y(n15) );
  AND2X2 U16 ( .A(n1155), .B(en), .Y(n16) );
  AND2X2 U17 ( .A(n519), .B(en), .Y(n17) );
  AND2X2 U18 ( .A(n678), .B(en), .Y(n18) );
  AND2X4 U19 ( .A(n25), .B(n26), .Y(temporary_overflow) );
  NAND2X1 U20 ( .A(output_p1_times_a1_mul_componentxinput_B_inverted_17_), 
        .B(n363), .Y(n20) );
  NAND2X1 U21 ( .A(input_p1_times_b1_mul_componentxinput_B_inverted_17_), 
        .B(n336), .Y(n21) );
  NAND2X1 U22 ( .A(input_p2_times_b2_mul_componentxinput_B_inverted_17_), 
        .B(n327), .Y(n22) );
  NAND2X1 U23 ( .A(output_p2_times_a2_mul_componentxinput_B_inverted_17_), 
        .B(n354), .Y(n23) );
  NAND2X1 U24 ( .A(input_times_b0_mul_componentxinput_B_inverted_17_), 
        .B(n345), .Y(n24) );
  NAND2X1 U25 ( .A(output_contracterxn1), .B(output_contracterxn2), .Y(n25) );
  NAND2X1 U26 ( .A(n27), .B(n28), .Y(n26) );
  INVX1 U27 ( .A(output_contracterxn4), .Y(n27) );
  INVX1 U28 ( .A(output_contracterxn3), .Y(n28) );
  XNOR2X4 U29 ( .A(n79), .B(n4168), .Y(\output_signal[1] ) );
  INVXL U30 ( .A(\output_signal[1] ), .Y(n1226) );
  INVX1 U31 ( .A(n348), .Y(n343) );
  INVX1 U32 ( .A(n342), .Y(n340) );
  INVX1 U33 ( .A(n333), .Y(n331) );
  INVX1 U34 ( .A(n324), .Y(n322) );
  INVX1 U35 ( .A(n360), .Y(n358) );
  INVX1 U36 ( .A(n351), .Y(n349) );
  INVX1 U37 ( .A(en), .Y(n370) );
  INVX1 U38 ( .A(en), .Y(n369) );
  INVX1 U39 ( .A(en), .Y(n372) );
  INVX1 U40 ( .A(en), .Y(n371) );
  INVX1 U41 ( .A(en), .Y(n367) );
  NOR2BX1 U42 ( .AN(n3817), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_15), .Y(n3816) );
  NAND2BX1 U43 ( .AN(output_p1_times_a1_mul_componentxunsigned_output_16), 
        .B(n3816), .Y(n3815) );
  INVX1 U44 ( .A(output_p1_times_a1_mul_componentxunsigned_output_9), .Y(n462)
         );
  NOR2BX1 U45 ( .AN(n3721), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_15), .Y(n3720) );
  NOR2BX1 U46 ( .AN(n3673), 
        .B(input_times_b0_mul_componentxunsigned_output_15), .Y(n3672) );
  NAND2BX1 U47 ( .AN(input_p1_times_b1_mul_componentxunsigned_output_16), 
        .B(n3720), .Y(n3719) );
  NAND2BX1 U48 ( .AN(input_p2_times_b2_mul_componentxunsigned_output_16), 
        .B(n3768), .Y(n3767) );
  NAND2BX1 U49 ( .AN(output_p2_times_a2_mul_componentxunsigned_output_16), 
        .B(n3864), .Y(n3863) );
  NAND2BX1 U50 ( .AN(input_times_b0_mul_componentxunsigned_output_16), 
        .B(n3672), .Y(n3671) );
  NOR2BX1 U51 ( .AN(n3769), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_15), .Y(n3768) );
  NOR2BX1 U52 ( .AN(n3865), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_15), .Y(n3864) );
  INVX1 U53 ( .A(input_p1_times_b1_mul_componentxunsigned_output_9), .Y(n939)
         );
  INVX1 U54 ( .A(input_p2_times_b2_mul_componentxunsigned_output_9), .Y(n1098)
         );
  INVX1 U55 ( .A(output_p2_times_a2_mul_componentxunsigned_output_9), .Y(n621)
         );
  INVX1 U56 ( .A(input_times_b0_mul_componentxunsigned_output_9), .Y(n780) );
  NOR3X1 U57 ( .A(output_p1_times_a1_mul_componentxunsigned_output_13), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_14), .C(n3818), 
        .Y(n3817) );
  XOR2X1 U58 ( .A(n2360), .B(n2361), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_14) );
  XOR2X1 U59 ( .A(n2356), .B(n2357), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_16) );
  XOR2X1 U60 ( .A(n2362), .B(n2363), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_13) );
  XOR2X1 U61 ( .A(n2349), .B(n2350), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_9) );
  XOR2X1 U62 ( .A(n2366), .B(n2367), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_11) );
  XOR2X1 U63 ( .A(n2358), .B(n2359), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_15) );
  XOR2X1 U64 ( .A(n2351), .B(n2352), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_8) );
  XOR2X1 U65 ( .A(n2364), .B(n2365), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_12) );
  XOR2X1 U66 ( .A(n2368), .B(n2369), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_10) );
  XOR2X1 U67 ( .A(n2316), .B(n2317), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_15) );
  XOR2X1 U68 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn518), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn519), 
        .Y(input_times_b0_mul_componentxunsigned_output_15) );
  XOR2X1 U69 ( .A(n2314), .B(n2315), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_16) );
  XOR2X1 U70 ( .A(n2335), .B(n2336), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_16) );
  XOR2X1 U71 ( .A(n2377), .B(n2378), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_16) );
  XOR2X1 U72 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn496), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn497), 
        .Y(input_times_b0_mul_componentxunsigned_output_16) );
  NOR3X1 U73 ( .A(input_p1_times_b1_mul_componentxunsigned_output_13), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_14), .C(n3722), 
        .Y(n3721) );
  NOR3X1 U74 ( .A(input_p2_times_b2_mul_componentxunsigned_output_13), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_14), .C(n3770), 
        .Y(n3769) );
  NOR3X1 U75 ( .A(output_p2_times_a2_mul_componentxunsigned_output_13), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_14), .C(n3866), 
        .Y(n3865) );
  NOR3X1 U76 ( .A(input_times_b0_mul_componentxunsigned_output_13), 
        .B(input_times_b0_mul_componentxunsigned_output_14), .C(n3674), 
        .Y(n3673) );
  XOR2X1 U77 ( .A(n2320), .B(n2321), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_13) );
  XOR2X1 U78 ( .A(n2341), .B(n2342), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_13) );
  XOR2X1 U79 ( .A(n2383), .B(n2384), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_13) );
  XOR2X1 U80 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn562), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn563), 
        .Y(input_times_b0_mul_componentxunsigned_output_13) );
  XOR2X1 U81 ( .A(n2307), .B(n2308), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_9) );
  XOR2X1 U82 ( .A(n2328), .B(n2329), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_9) );
  XOR2X1 U83 ( .A(n2370), .B(n2371), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_9) );
  XOR2X1 U84 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn2), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn3), 
        .Y(input_times_b0_mul_componentxunsigned_output_9) );
  XOR2X1 U85 ( .A(n2324), .B(n2325), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_11) );
  XOR2X1 U86 ( .A(n2345), .B(n2346), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_11) );
  XOR2X1 U87 ( .A(n2387), .B(n2388), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_11) );
  XOR2X1 U88 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn606), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn607), 
        .Y(input_times_b0_mul_componentxunsigned_output_11) );
  XOR2X1 U89 ( .A(n2337), .B(n2338), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_15) );
  XOR2X1 U90 ( .A(n2379), .B(n2380), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_15) );
  XOR2X1 U91 ( .A(n2309), .B(n2310), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_8) );
  XOR2X1 U92 ( .A(n2318), .B(n2319), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_14) );
  XOR2X1 U93 ( .A(n2330), .B(n2331), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_8) );
  XOR2X1 U94 ( .A(n2339), .B(n2340), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_14) );
  XOR2X1 U95 ( .A(n2372), .B(n2373), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_8) );
  XOR2X1 U96 ( .A(n2381), .B(n2382), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_14) );
  XOR2X1 U97 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn24), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn25), 
        .Y(input_times_b0_mul_componentxunsigned_output_8) );
  XOR2X1 U98 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn540), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn541), 
        .Y(input_times_b0_mul_componentxunsigned_output_14) );
  XOR2X1 U99 ( .A(n2322), .B(n2323), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_12) );
  XOR2X1 U100 ( .A(n2343), .B(n2344), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_12) );
  XOR2X1 U101 ( .A(n2385), .B(n2386), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_12) );
  XOR2X1 U102 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn584), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn585), 
        .Y(input_times_b0_mul_componentxunsigned_output_12) );
  XOR2X1 U103 ( .A(n2326), .B(n2327), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_10) );
  XOR2X1 U104 ( .A(n2347), .B(n2348), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_10) );
  XOR2X1 U105 ( .A(n2389), .B(n2390), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_10) );
  XOR2X1 U106 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn628), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn629), 
        .Y(input_times_b0_mul_componentxunsigned_output_10) );
  AOI22X1 U107 ( .A0(output_p1_times_a1_mul_componentxUMxsecond_vector[9]), 
        .A1(output_p1_times_a1_mul_componentxUMxfirst_vector[9]), .B0(n2349), 
        .B1(n2350), .Y(n2369) );
  AOI22X1 U108 ( .A0(output_p1_times_a1_mul_componentxUMxsecond_vector[11]), 
        .A1(output_p1_times_a1_mul_componentxUMxfirst_vector[11]), .B0(n2366), 
        .B1(n2367), .Y(n2365) );
  AOI22X1 U109 ( .A0(output_p1_times_a1_mul_componentxUMxsecond_vector[13]), 
        .A1(output_p1_times_a1_mul_componentxUMxfirst_vector[13]), .B0(n2362), 
        .B1(n2363), .Y(n2361) );
  AOI22X1 U110 ( .A0(output_p1_times_a1_mul_componentxUMxsecond_vector[15]), 
        .A1(output_p1_times_a1_mul_componentxUMxfirst_vector[15]), .B0(n2358), 
        .B1(n2359), .Y(n2357) );
  OAI2BB2X1 U111 ( .B0(n2365), .B1(n2364), 
        .A0N(output_p1_times_a1_mul_componentxUMxsecond_vector[12]), 
        .A1N(output_p1_times_a1_mul_componentxUMxfirst_vector[12]), .Y(n2362)
         );
  OAI2BB2X1 U112 ( .B0(n2361), .B1(n2360), 
        .A0N(output_p1_times_a1_mul_componentxUMxsecond_vector[14]), 
        .A1N(output_p1_times_a1_mul_componentxUMxfirst_vector[14]), .Y(n2358)
         );
  OAI2BB2X1 U113 ( .B0(n2369), .B1(n2368), 
        .A0N(output_p1_times_a1_mul_componentxUMxsecond_vector[10]), 
        .A1N(output_p1_times_a1_mul_componentxUMxfirst_vector[10]), .Y(n2366)
         );
  OAI2BB2X1 U114 ( .B0(n2352), .B1(n2351), 
        .A0N(output_p1_times_a1_mul_componentxUMxsecond_vector[8]), 
        .A1N(output_p1_times_a1_mul_componentxUMxfirst_vector[8]), .Y(n2349)
         );
  OAI2BB2X1 U115 ( .B0(n2357), .B1(n2356), 
        .A0N(output_p1_times_a1_mul_componentxUMxsecond_vector[16]), 
        .A1N(n407), .Y(n2354) );
  XNOR2X1 U116 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[8]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[8]), .Y(n2351) );
  XOR2X1 U117 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[7]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[7]), .Y(n2353) );
  NAND2X1 U118 ( .A(output_p1_times_a1_mul_componentxUMxsecond_vector[7]), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[7]), .Y(n2352) );
  XOR2X1 U119 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .B(n3320), .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[15])
         );
  XOR2X1 U120 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[9]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[9]), .Y(n2350) );
  XOR2X1 U121 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[11]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[11]), .Y(n2367)
         );
  XOR2X1 U122 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[13]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[13]), .Y(n2363)
         );
  XOR2X1 U123 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[15]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[15]), .Y(n2359)
         );
  OR3XL U124 ( .A(output_p1_times_a1_mul_componentxunsigned_output_11), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_12), .C(n3820), 
        .Y(n3818) );
  XNOR2X1 U125 ( .A(n407), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[16]), .Y(n2356)
         );
  XNOR2X1 U126 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[10]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[10]), .Y(n2368)
         );
  XNOR2X1 U127 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[12]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[12]), .Y(n2364)
         );
  XNOR2X1 U128 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[14]), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[14]), .Y(n2360)
         );
  XOR2X1 U129 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .B(n3322), .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[16])
         );
  AOI22X1 U130 ( .A0(input_p1_times_b1_mul_componentxUMxsecond_vector[13]), 
        .A1(input_p1_times_b1_mul_componentxUMxfirst_vector[13]), .B0(n2320), 
        .B1(n2321), .Y(n2319) );
  AOI22X1 U131 ( .A0(input_times_b0_mul_componentxUMxsecond_vector[13]), 
        .A1(input_times_b0_mul_componentxUMxfirst_vector[13]), 
        .B0(input_times_b0_mul_componentxUMxAdder_finalxn562), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn563), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn541) );
  AOI22X1 U132 ( .A0(input_p1_times_b1_mul_componentxUMxsecond_vector[15]), 
        .A1(input_p1_times_b1_mul_componentxUMxfirst_vector[15]), .B0(n2316), 
        .B1(n2317), .Y(n2315) );
  AOI22X1 U133 ( .A0(input_p2_times_b2_mul_componentxUMxsecond_vector[15]), 
        .A1(input_p2_times_b2_mul_componentxUMxfirst_vector[15]), .B0(n2337), 
        .B1(n2338), .Y(n2336) );
  AOI22X1 U134 ( .A0(output_p2_times_a2_mul_componentxUMxsecond_vector[15]), 
        .A1(output_p2_times_a2_mul_componentxUMxfirst_vector[15]), .B0(n2379), 
        .B1(n2380), .Y(n2378) );
  AOI22X1 U135 ( .A0(input_times_b0_mul_componentxUMxsecond_vector[15]), 
        .A1(input_times_b0_mul_componentxUMxfirst_vector[15]), 
        .B0(input_times_b0_mul_componentxUMxAdder_finalxn518), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn519), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn497) );
  OAI2BB2X1 U136 ( .B0(n2319), .B1(n2318), 
        .A0N(input_p1_times_b1_mul_componentxUMxsecond_vector[14]), 
        .A1N(input_p1_times_b1_mul_componentxUMxfirst_vector[14]), .Y(n2316)
         );
  OAI2BB2X1 U137 ( .B0(input_times_b0_mul_componentxUMxAdder_finalxn541), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn540), 
        .A0N(input_times_b0_mul_componentxUMxsecond_vector[14]), 
        .A1N(input_times_b0_mul_componentxUMxfirst_vector[14]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn518) );
  OAI2BB2X1 U138 ( .B0(n2315), .B1(n2314), 
        .A0N(input_p1_times_b1_mul_componentxUMxsecond_vector[16]), .A1N(n883), 
        .Y(n2312) );
  OAI2BB2X1 U139 ( .B0(n2336), .B1(n2335), 
        .A0N(input_p2_times_b2_mul_componentxUMxsecond_vector[16]), 
        .A1N(n1042), .Y(n2333) );
  OAI2BB2X1 U140 ( .B0(n2378), .B1(n2377), 
        .A0N(output_p2_times_a2_mul_componentxUMxsecond_vector[16]), 
        .A1N(n565), .Y(n2375) );
  OAI2BB2X1 U141 ( .B0(input_times_b0_mul_componentxUMxAdder_finalxn497), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn496), 
        .A0N(input_times_b0_mul_componentxUMxsecond_vector[16]), .A1N(n724), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn474) );
  XOR2X1 U142 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .B(n2852), .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[15]) );
  XOR2X1 U143 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .B(n3086), .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[15]) );
  XOR2X1 U144 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .B(n3554), .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[15])
         );
  XOR2X1 U145 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .B(n2618), .Y(input_times_b0_mul_componentxUMxsecond_vector[15]) );
  XOR2X1 U146 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[13]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[13]), .Y(n2321) );
  XOR2X1 U147 ( .A(input_times_b0_mul_componentxUMxfirst_vector[13]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[13]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn563) );
  XOR2X1 U148 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[15]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[15]), .Y(n2317) );
  XOR2X1 U149 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[15]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[15]), .Y(n2338) );
  XOR2X1 U150 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[15]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[15]), .Y(n2380)
         );
  XOR2X1 U151 ( .A(input_times_b0_mul_componentxUMxfirst_vector[15]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[15]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn519) );
  XNOR2X1 U152 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[14]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[14]), .Y(n2318) );
  XNOR2X1 U153 ( .A(input_times_b0_mul_componentxUMxfirst_vector[14]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[14]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn540) );
  AOI22X1 U154 ( .A0(input_p1_times_b1_mul_componentxUMxsecond_vector[9]), 
        .A1(input_p1_times_b1_mul_componentxUMxfirst_vector[9]), .B0(n2307), 
        .B1(n2308), .Y(n2327) );
  AOI22X1 U155 ( .A0(input_p2_times_b2_mul_componentxUMxsecond_vector[9]), 
        .A1(input_p2_times_b2_mul_componentxUMxfirst_vector[9]), .B0(n2328), 
        .B1(n2329), .Y(n2348) );
  AOI22X1 U156 ( .A0(output_p2_times_a2_mul_componentxUMxsecond_vector[9]), 
        .A1(output_p2_times_a2_mul_componentxUMxfirst_vector[9]), .B0(n2370), 
        .B1(n2371), .Y(n2390) );
  AOI22X1 U157 ( .A0(input_times_b0_mul_componentxUMxsecond_vector[9]), 
        .A1(input_times_b0_mul_componentxUMxfirst_vector[9]), 
        .B0(input_times_b0_mul_componentxUMxAdder_finalxn2), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn3), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn629) );
  AOI22X1 U158 ( .A0(input_p1_times_b1_mul_componentxUMxsecond_vector[11]), 
        .A1(input_p1_times_b1_mul_componentxUMxfirst_vector[11]), .B0(n2324), 
        .B1(n2325), .Y(n2323) );
  AOI22X1 U159 ( .A0(input_p2_times_b2_mul_componentxUMxsecond_vector[11]), 
        .A1(input_p2_times_b2_mul_componentxUMxfirst_vector[11]), .B0(n2345), 
        .B1(n2346), .Y(n2344) );
  AOI22X1 U160 ( .A0(output_p2_times_a2_mul_componentxUMxsecond_vector[11]), 
        .A1(output_p2_times_a2_mul_componentxUMxfirst_vector[11]), .B0(n2387), 
        .B1(n2388), .Y(n2386) );
  AOI22X1 U161 ( .A0(input_times_b0_mul_componentxUMxsecond_vector[11]), 
        .A1(input_times_b0_mul_componentxUMxfirst_vector[11]), 
        .B0(input_times_b0_mul_componentxUMxAdder_finalxn606), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn607), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn585) );
  AOI22X1 U162 ( .A0(input_p2_times_b2_mul_componentxUMxsecond_vector[13]), 
        .A1(input_p2_times_b2_mul_componentxUMxfirst_vector[13]), .B0(n2341), 
        .B1(n2342), .Y(n2340) );
  AOI22X1 U163 ( .A0(output_p2_times_a2_mul_componentxUMxsecond_vector[13]), 
        .A1(output_p2_times_a2_mul_componentxUMxfirst_vector[13]), .B0(n2383), 
        .B1(n2384), .Y(n2382) );
  OAI2BB2X1 U164 ( .B0(n2323), .B1(n2322), 
        .A0N(input_p1_times_b1_mul_componentxUMxsecond_vector[12]), 
        .A1N(input_p1_times_b1_mul_componentxUMxfirst_vector[12]), .Y(n2320)
         );
  OAI2BB2X1 U165 ( .B0(n2344), .B1(n2343), 
        .A0N(input_p2_times_b2_mul_componentxUMxsecond_vector[12]), 
        .A1N(input_p2_times_b2_mul_componentxUMxfirst_vector[12]), .Y(n2341)
         );
  OAI2BB2X1 U166 ( .B0(n2386), .B1(n2385), 
        .A0N(output_p2_times_a2_mul_componentxUMxsecond_vector[12]), 
        .A1N(output_p2_times_a2_mul_componentxUMxfirst_vector[12]), .Y(n2383)
         );
  OAI2BB2X1 U167 ( .B0(input_times_b0_mul_componentxUMxAdder_finalxn585), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn584), 
        .A0N(input_times_b0_mul_componentxUMxsecond_vector[12]), 
        .A1N(input_times_b0_mul_componentxUMxfirst_vector[12]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn562) );
  OAI2BB2X1 U168 ( .B0(n2340), .B1(n2339), 
        .A0N(input_p2_times_b2_mul_componentxUMxsecond_vector[14]), 
        .A1N(input_p2_times_b2_mul_componentxUMxfirst_vector[14]), .Y(n2337)
         );
  OAI2BB2X1 U169 ( .B0(n2382), .B1(n2381), 
        .A0N(output_p2_times_a2_mul_componentxUMxsecond_vector[14]), 
        .A1N(output_p2_times_a2_mul_componentxUMxfirst_vector[14]), .Y(n2379)
         );
  OAI2BB2X1 U170 ( .B0(n2327), .B1(n2326), 
        .A0N(input_p1_times_b1_mul_componentxUMxsecond_vector[10]), 
        .A1N(input_p1_times_b1_mul_componentxUMxfirst_vector[10]), .Y(n2324)
         );
  OAI2BB2X1 U171 ( .B0(n2348), .B1(n2347), 
        .A0N(input_p2_times_b2_mul_componentxUMxsecond_vector[10]), 
        .A1N(input_p2_times_b2_mul_componentxUMxfirst_vector[10]), .Y(n2345)
         );
  OAI2BB2X1 U172 ( .B0(n2390), .B1(n2389), 
        .A0N(output_p2_times_a2_mul_componentxUMxsecond_vector[10]), 
        .A1N(output_p2_times_a2_mul_componentxUMxfirst_vector[10]), .Y(n2387)
         );
  OAI2BB2X1 U173 ( .B0(input_times_b0_mul_componentxUMxAdder_finalxn629), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn628), 
        .A0N(input_times_b0_mul_componentxUMxsecond_vector[10]), 
        .A1N(input_times_b0_mul_componentxUMxfirst_vector[10]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn606) );
  OAI2BB2X1 U174 ( .B0(n2310), .B1(n2309), 
        .A0N(input_p1_times_b1_mul_componentxUMxsecond_vector[8]), 
        .A1N(input_p1_times_b1_mul_componentxUMxfirst_vector[8]), .Y(n2307) );
  OAI2BB2X1 U175 ( .B0(n2331), .B1(n2330), 
        .A0N(input_p2_times_b2_mul_componentxUMxsecond_vector[8]), 
        .A1N(input_p2_times_b2_mul_componentxUMxfirst_vector[8]), .Y(n2328) );
  OAI2BB2X1 U176 ( .B0(n2373), .B1(n2372), 
        .A0N(output_p2_times_a2_mul_componentxUMxsecond_vector[8]), 
        .A1N(output_p2_times_a2_mul_componentxUMxfirst_vector[8]), .Y(n2370)
         );
  OAI2BB2X1 U177 ( .B0(input_times_b0_mul_componentxUMxAdder_finalxn25), 
        .B1(input_times_b0_mul_componentxUMxAdder_finalxn24), 
        .A0N(input_times_b0_mul_componentxUMxsecond_vector[8]), 
        .A1N(input_times_b0_mul_componentxUMxfirst_vector[8]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn2) );
  NAND2X1 U178 ( .A(input_p1_times_b1_mul_componentxUMxsecond_vector[7]), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[7]), .Y(n2310) );
  NAND2X1 U179 ( .A(input_p2_times_b2_mul_componentxUMxsecond_vector[7]), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[7]), .Y(n2331) );
  NAND2X1 U180 ( .A(output_p2_times_a2_mul_componentxUMxsecond_vector[7]), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[7]), .Y(n2373) );
  NAND2X1 U181 ( .A(input_times_b0_mul_componentxUMxsecond_vector[7]), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[7]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn25) );
  XOR2X1 U182 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[9]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[9]), .Y(n2308) );
  XOR2X1 U183 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[9]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[9]), .Y(n2329) );
  XOR2X1 U184 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[9]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[9]), .Y(n2371) );
  XOR2X1 U185 ( .A(input_times_b0_mul_componentxUMxfirst_vector[9]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[9]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn3) );
  XOR2X1 U186 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[11]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[11]), .Y(n2325) );
  XOR2X1 U187 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[11]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[11]), .Y(n2346) );
  XOR2X1 U188 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[11]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[11]), .Y(n2388)
         );
  XOR2X1 U189 ( .A(input_times_b0_mul_componentxUMxfirst_vector[11]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[11]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn607) );
  XOR2X1 U190 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[13]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[13]), .Y(n2342) );
  XOR2X1 U191 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[13]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[13]), .Y(n2384)
         );
  OR3XL U192 ( .A(input_p1_times_b1_mul_componentxunsigned_output_11), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_12), .C(n3724), 
        .Y(n3722) );
  OR3XL U193 ( .A(input_p2_times_b2_mul_componentxunsigned_output_11), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_12), .C(n3772), 
        .Y(n3770) );
  OR3XL U194 ( .A(output_p2_times_a2_mul_componentxunsigned_output_11), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_12), .C(n3868), 
        .Y(n3866) );
  OR3XL U195 ( .A(input_times_b0_mul_componentxunsigned_output_11), 
        .B(input_times_b0_mul_componentxunsigned_output_12), .C(n3676), 
        .Y(n3674) );
  XNOR2X1 U196 ( .A(n883), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[16]), .Y(n2314) );
  XNOR2X1 U197 ( .A(n1042), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[16]), .Y(n2335) );
  XNOR2X1 U198 ( .A(n565), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[16]), .Y(n2377)
         );
  XNOR2X1 U199 ( .A(n724), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[16]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn496) );
  XNOR2X1 U200 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[8]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[8]), .Y(n2309) );
  XNOR2X1 U201 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[8]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[8]), .Y(n2330) );
  XNOR2X1 U202 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[8]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[8]), .Y(n2372) );
  XNOR2X1 U203 ( .A(input_times_b0_mul_componentxUMxfirst_vector[8]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[8]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn24) );
  XNOR2X1 U204 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[10]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[10]), .Y(n2326) );
  XNOR2X1 U205 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[10]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[10]), .Y(n2347) );
  XNOR2X1 U206 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[10]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[10]), .Y(n2389)
         );
  XNOR2X1 U207 ( .A(input_times_b0_mul_componentxUMxfirst_vector[10]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[10]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn628) );
  XNOR2X1 U208 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[12]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[12]), .Y(n2322) );
  XNOR2X1 U209 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[12]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[12]), .Y(n2343) );
  XNOR2X1 U210 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[12]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[12]), .Y(n2385)
         );
  XNOR2X1 U211 ( .A(input_times_b0_mul_componentxUMxfirst_vector[12]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[12]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn584) );
  XNOR2X1 U212 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[14]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[14]), .Y(n2339) );
  XNOR2X1 U213 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[14]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[14]), .Y(n2381)
         );
  XOR2X1 U214 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .B(n2854), .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[16]) );
  XOR2X1 U215 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .B(n3088), .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[16]) );
  XOR2X1 U216 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .B(n3556), .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[16])
         );
  XOR2X1 U217 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .B(n2620), .Y(input_times_b0_mul_componentxUMxsecond_vector[16]) );
  XOR2X1 U218 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[7]), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[7]), .Y(n2311) );
  XOR2X1 U219 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[7]), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[7]), .Y(n2332) );
  XOR2X1 U220 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[7]), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[7]), .Y(n2374) );
  XOR2X1 U221 ( .A(input_times_b0_mul_componentxUMxfirst_vector[7]), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[7]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn47) );
  XOR2X1 U222 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[8]) );
  NAND3BX1 U223 ( .AN(output_p1_times_a1_mul_componentxunsigned_output_10), 
        .B(n462), .C(n3807), .Y(n3820) );
  XOR2X1 U224 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[6]) );
  XOR2X1 U225 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[9]) );
  XOR2X1 U226 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n452), .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[11]) );
  XOR2X1 U227 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n431), .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[13]) );
  XOR2X1 U228 ( .A(n429), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .Y(n3313) );
  XOR2X1 U229 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B(n416), .Y(n3320) );
  XOR2X1 U230 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B(n414), .Y(n3322) );
  XOR2X1 U231 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[7]) );
  XOR2X1 U232 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[10]) );
  XOR2X1 U233 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n440), .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[12]) );
  XOR2X1 U234 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n422), .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[14]) );
  XOR2X1 U235 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .B(n3315), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128220800_128221024_128221136)
         );
  AND2X2 U236 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[9]) );
  AND2X2 U237 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[11]) );
  AND2X2 U238 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n440), .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[13]) );
  AND2X2 U239 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[7]) );
  XOR2X1 U240 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .B(n3305), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128125248_128219960_128220240)
         );
  XOR2X1 U241 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .B(n3307), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128125584_128220184_128220408)
         );
  XOR2X1 U242 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .B(n3309), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128125920_128220352_128220576)
         );
  XOR2X1 U243 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .B(n3311), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128126256_128220520_128220744)
         );
  XOR2X1 U244 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128126480_128126592), 
        .B(n3313), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128220688_128220856_128220968)
         );
  AND2X2 U245 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[8]) );
  AND2X2 U246 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[10]) );
  AND2X2 U247 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n452), .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[12]) );
  AND2X2 U248 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n431), .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[14]) );
  INVX1 U249 ( .A(n3314), .Y(n416) );
  AOI22X1 U250 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .A1(n429), .B0(n3313), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer4_128126480_128126592), 
        .Y(n3314) );
  INVX1 U251 ( .A(n3321), .Y(n407) );
  AOI22X1 U252 ( .A0(n416), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B0(n3320), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .Y(n3321) );
  AOI22X1 U253 ( .A0(n414), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B0(n3322), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .Y(n3323) );
  XOR2X1 U254 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .B(n3317), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128315464_128315632_128315800)
         );
  AND2X2 U255 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n422), .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[15]) );
  INVX1 U256 ( .A(n2846), .Y(n892) );
  AOI22X1 U257 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .A1(n905), .B0(n2845), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer4_128126480_128126592), 
        .Y(n2846) );
  INVX1 U258 ( .A(n2612), .Y(n733) );
  AOI22X1 U259 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .A1(n746), .B0(n2611), 
        .B1(input_times_b0_mul_componentxUMxsum_layer4_128126480_128126592), 
        .Y(n2612) );
  XOR2X1 U260 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n907), .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[13]) );
  XOR2X1 U261 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n748), .Y(input_times_b0_mul_componentxUMxsecond_vector[13]) );
  XOR2X1 U262 ( .A(n905), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .Y(n2845) );
  XOR2X1 U263 ( .A(n1064), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .Y(n3079) );
  XOR2X1 U264 ( .A(n587), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .Y(n3547) );
  XOR2X1 U265 ( .A(n746), 
        .B(input_times_b0_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .Y(n2611) );
  XOR2X1 U266 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B(n892), .Y(n2852) );
  XOR2X1 U267 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B(n1051), .Y(n3086) );
  XOR2X1 U268 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B(n574), .Y(n3554) );
  XOR2X1 U269 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B(n733), .Y(n2618) );
  XOR2X1 U270 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n898), .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[14]) );
  XOR2X1 U271 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n739), .Y(input_times_b0_mul_componentxUMxsecond_vector[14]) );
  XOR2X1 U272 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .B(n2843), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128126256_128220520_128220744)
         );
  XOR2X1 U273 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .B(n2609), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128126256_128220520_128220744)
         );
  XOR2X1 U274 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128126480_128126592), 
        .B(n2845), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128220688_128220856_128220968)
         );
  XOR2X1 U275 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128126480_128126592), 
        .B(n2611), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128220688_128220856_128220968)
         );
  INVX1 U276 ( .A(n3080), .Y(n1051) );
  AOI22X1 U277 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .A1(n1064), .B0(n3079), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer4_128126480_128126592), 
        .Y(n3080) );
  INVX1 U278 ( .A(n3548), .Y(n574) );
  AOI22X1 U279 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer4_128262496_128126088_128126312), 
        .A1(n587), .B0(n3547), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer4_128126480_128126592), 
        .Y(n3548) );
  AOI22X1 U280 ( .A0(n890), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B0(n2854), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .Y(n2855) );
  AOI22X1 U281 ( .A0(n1049), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B0(n3088), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .Y(n3089) );
  AOI22X1 U282 ( .A0(n572), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B0(n3556), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .Y(n3557) );
  AOI22X1 U283 ( .A0(n731), 
        .A1(input_times_b0_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B0(n2620), 
        .B1(input_times_b0_mul_componentxUMxsum_layer5_128315464_128315632_128315800), 
        .Y(n2621) );
  NAND3BX1 U284 ( .AN(input_p1_times_b1_mul_componentxunsigned_output_10), 
        .B(n939), .C(n3711), .Y(n3724) );
  NAND3BX1 U285 ( .AN(input_p2_times_b2_mul_componentxunsigned_output_10), 
        .B(n1098), .C(n3759), .Y(n3772) );
  NAND3BX1 U286 ( .AN(output_p2_times_a2_mul_componentxunsigned_output_10), 
        .B(n621), .C(n3855), .Y(n3868) );
  NAND3BX1 U287 ( .AN(input_times_b0_mul_componentxunsigned_output_10), 
        .B(n780), .C(n3663), .Y(n3676) );
  XOR2X1 U288 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[9]) );
  XOR2X1 U289 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[9]) );
  XOR2X1 U290 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[9]) );
  XOR2X1 U291 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(input_times_b0_mul_componentxUMxsecond_vector[9]) );
  XOR2X1 U292 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n929), .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[11]) );
  XOR2X1 U293 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n1088), .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[11]) );
  XOR2X1 U294 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n611), .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[11]) );
  XOR2X1 U295 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n770), .Y(input_times_b0_mul_componentxUMxsecond_vector[11]) );
  XOR2X1 U296 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n1066), .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[13]) );
  XOR2X1 U297 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n589), .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[13]) );
  XOR2X1 U298 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B(n890), .Y(n2854) );
  XOR2X1 U299 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B(n1049), .Y(n3088) );
  XOR2X1 U300 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B(n572), .Y(n3556) );
  XOR2X1 U301 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128237920_128238088), 
        .B(n731), .Y(n2620) );
  XOR2X1 U302 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[7]) );
  XOR2X1 U303 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[7]) );
  XOR2X1 U304 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[7]) );
  XOR2X1 U305 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(input_times_b0_mul_componentxUMxsecond_vector[7]) );
  XOR2X1 U306 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[8]) );
  XOR2X1 U307 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[8]) );
  XOR2X1 U308 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[8]) );
  XOR2X1 U309 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(input_times_b0_mul_componentxUMxsecond_vector[8]) );
  XOR2X1 U310 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[10]) );
  XOR2X1 U311 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[10]) );
  XOR2X1 U312 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[10]) );
  XOR2X1 U313 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(input_times_b0_mul_componentxUMxsecond_vector[10]) );
  XOR2X1 U314 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n916), .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[12]) );
  XOR2X1 U315 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n1075), .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[12]) );
  XOR2X1 U316 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n598), .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[12]) );
  XOR2X1 U317 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n757), .Y(input_times_b0_mul_componentxUMxsecond_vector[12]) );
  XOR2X1 U318 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n1057), .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[14]) );
  XOR2X1 U319 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n580), .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[14]) );
  XOR2X1 U320 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .B(n2847), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128220800_128221024_128221136)
         );
  XOR2X1 U321 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .B(n3081), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128220800_128221024_128221136)
         );
  XOR2X1 U322 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .B(n3549), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128220800_128221024_128221136)
         );
  XOR2X1 U323 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .B(n2613), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128220800_128221024_128221136)
         );
  XOR2X1 U324 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .B(n2849), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128315464_128315632_128315800)
         );
  XOR2X1 U325 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .B(n3083), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128315464_128315632_128315800)
         );
  XOR2X1 U326 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .B(n3551), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128315464_128315632_128315800)
         );
  XOR2X1 U327 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .B(n2615), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128315464_128315632_128315800)
         );
  AND2X2 U328 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[9]) );
  AND2X2 U329 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[9]) );
  AND2X2 U330 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[9]) );
  AND2X2 U331 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128219624_128219848), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219456_128219680), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[9]) );
  AND2X2 U332 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[11]) );
  AND2X2 U333 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[11]) );
  AND2X2 U334 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[11]) );
  AND2X2 U335 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128125248_128219960_128220240), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219792_128220016), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[11]) );
  AND2X2 U336 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n916), .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[13]) );
  AND2X2 U337 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n1075), .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[13]) );
  AND2X2 U338 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n598), .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[13]) );
  AND2X2 U339 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128125920_128220352_128220576), 
        .B(n757), .Y(input_times_b0_mul_componentxUMxfirst_vector[13]) );
  AND2X2 U340 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n898), .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[15]) );
  AND2X2 U341 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n1057), .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[15]) );
  AND2X2 U342 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n580), .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[15]) );
  AND2X2 U343 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128220688_128220856_128220968), 
        .B(n739), .Y(input_times_b0_mul_componentxUMxfirst_vector[15]) );
  AND2X2 U344 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[7]) );
  AND2X2 U345 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[7]) );
  XOR2X1 U346 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .B(n2837), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128125248_128219960_128220240)
         );
  XOR2X1 U347 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .B(n3071), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128125248_128219960_128220240)
         );
  XOR2X1 U348 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .B(n3539), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128125248_128219960_128220240)
         );
  XOR2X1 U349 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .B(n2603), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128125248_128219960_128220240)
         );
  XOR2X1 U350 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .B(n2839), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128125584_128220184_128220408)
         );
  XOR2X1 U351 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .B(n3073), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128125584_128220184_128220408)
         );
  XOR2X1 U352 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .B(n3541), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128125584_128220184_128220408)
         );
  XOR2X1 U353 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .B(n2605), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128125584_128220184_128220408)
         );
  XOR2X1 U354 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .B(n2841), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128125920_128220352_128220576)
         );
  XOR2X1 U355 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .B(n3075), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128125920_128220352_128220576)
         );
  XOR2X1 U356 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .B(n3543), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128125920_128220352_128220576)
         );
  XOR2X1 U357 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .B(n2607), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128125920_128220352_128220576)
         );
  XOR2X1 U358 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .B(n3077), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128126256_128220520_128220744)
         );
  XOR2X1 U359 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .B(n3545), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128126256_128220520_128220744)
         );
  XOR2X1 U360 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128126480_128126592), 
        .B(n3079), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128220688_128220856_128220968)
         );
  XOR2X1 U361 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128126480_128126592), 
        .B(n3547), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128220688_128220856_128220968)
         );
  AND2X2 U362 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[8]) );
  AND2X2 U363 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[8]) );
  AND2X2 U364 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[8]) );
  AND2X2 U365 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128219456_128219680), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219288_128219512), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[8]) );
  AND2X2 U366 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[10]) );
  AND2X2 U367 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[10]) );
  AND2X2 U368 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[10]) );
  AND2X2 U369 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128219792_128220016), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219624_128219848), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[10]) );
  AND2X2 U370 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n929), .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[12]) );
  AND2X2 U371 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n1088), .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[12]) );
  AND2X2 U372 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n611), .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[12]) );
  AND2X2 U373 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128125584_128220184_128220408), 
        .B(n770), .Y(input_times_b0_mul_componentxUMxfirst_vector[12]) );
  AND2X2 U374 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n907), .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[14]) );
  AND2X2 U375 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n1066), .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[14]) );
  AND2X2 U376 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n589), .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[14]) );
  AND2X2 U377 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128126256_128220520_128220744), 
        .B(n748), .Y(input_times_b0_mul_componentxUMxfirst_vector[14]) );
  INVX1 U378 ( .A(n2853), .Y(n883) );
  AOI22X1 U379 ( .A0(n892), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B0(n2852), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .Y(n2853) );
  INVX1 U380 ( .A(n3087), .Y(n1042) );
  AOI22X1 U381 ( .A0(n1051), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B0(n3086), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .Y(n3087) );
  INVX1 U382 ( .A(n3555), .Y(n565) );
  AOI22X1 U383 ( .A0(n574), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B0(n3554), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .Y(n3555) );
  INVX1 U384 ( .A(n2619), .Y(n724) );
  AOI22X1 U385 ( .A0(n733), 
        .A1(input_times_b0_mul_componentxUMxsum_layer4_128126816_128126928), 
        .B0(n2618), 
        .B1(input_times_b0_mul_componentxUMxsum_layer5_128220800_128221024_128221136), 
        .Y(n2619) );
  XOR2X1 U386 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[6]) );
  XOR2X1 U387 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[6]) );
  XOR2X1 U388 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[6]) );
  XOR2X1 U389 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(input_times_b0_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[6]) );
  AND2X2 U390 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[7]) );
  AND2X2 U391 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128219288_128219512), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219120_128219344), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[7]) );
  AND2X2 U392 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219456_128219680)
         );
  XOR2X1 U393 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .B(n3285), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128247456_128124464_128124688)
         );
  XOR2X1 U394 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .B(n3283), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128247120_128124240_128124520)
         );
  XOR2X1 U395 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n481), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128219624_128219848)
         );
  BUFX3 U396 ( .A(n398), .Y(n112) );
  BUFX3 U397 ( .A(n398), .Y(n111) );
  NOR3X1 U398 ( .A(\output_signal[7] ), .B(output_previous_1[8]), .C(n3777), 
        .Y(n3775) );
  NOR3X1 U399 ( .A(n2353), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_8), .C(n3809), 
        .Y(n3807) );
  NAND3BX1 U400 ( .AN(output_previous_1[10]), .B(n1210), .C(n3775), .Y(n3788)
         );
  INVX1 U401 ( .A(n3296), .Y(n429) );
  AOI22X1 U402 ( .A0(n430), .A1(n437), .B0(n3295), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .Y(n3296) );
  OR3XL U403 ( .A(\output_signal[5] ), .B(\output_signal[6] ), .C(n3779), 
        .Y(n3777) );
  XOR2X1 U404 ( .A(n421), .B(n3297), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128262496_128126088_128126312)
         );
  XOR2X1 U405 ( .A(n478), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .Y(n3287) );
  XOR2X1 U406 ( .A(n449), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .Y(n3293) );
  XOR2X1 U407 ( .A(n415), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .Y(n3315) );
  XOR2X1 U408 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B(n464), .Y(n3305) );
  XOR2X1 U409 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B(n460), .Y(n3307) );
  XOR2X1 U410 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B(n448), .Y(n3309) );
  XOR2X1 U411 ( .A(n437), .B(n430), .Y(n3295) );
  XOR2X1 U412 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B(n438), .Y(n3311) );
  XOR2X1 U413 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .B(n3289), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128124744_128124968_128125136)
         );
  XOR2X1 U414 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .B(n3291), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128125080_128125304_128125472)
         );
  XOR2X1 U415 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .B(n3293), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128125416_128125640_128125808)
         );
  XOR2X1 U416 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .B(n3295), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128125752_128125976_128126144)
         );
  AND2X2 U417 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219288_128219512)
         );
  AND2X2 U418 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219120_128219344)
         );
  AND2X2 U419 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n481), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219624_128219848)
         );
  AND2X2 U420 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n472), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer5_128219792_128220016)
         );
  XOR2X1 U421 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128219456_128219680)
         );
  XOR2X1 U422 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128219288_128219512)
         );
  XOR2X1 U423 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128247680_128247792), 
        .B(n3287), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128124632_128124800_128124912)
         );
  XOR2X1 U424 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n472), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128219792_128220016)
         );
  INVX1 U425 ( .A(n3288), .Y(n464) );
  AOI22X1 U426 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .A1(n478), .B0(n3287), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer3_128247680_128247792), 
        .Y(n3288) );
  INVX1 U427 ( .A(n3294), .Y(n438) );
  AOI22X1 U428 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .A1(n449), .B0(n3293), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .Y(n3294) );
  INVX1 U429 ( .A(n3316), .Y(n414) );
  AOI22X1 U430 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .A1(n415), .B0(n3315), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .Y(n3316) );
  INVX1 U431 ( .A(n3306), .Y(n452) );
  AOI22X1 U432 ( .A0(n464), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B0(n3305), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .Y(n3306) );
  INVX1 U433 ( .A(n3308), .Y(n440) );
  AOI22X1 U434 ( .A0(n460), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B0(n3307), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .Y(n3308) );
  INVX1 U435 ( .A(n3310), .Y(n431) );
  AOI22X1 U436 ( .A0(n448), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B0(n3309), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .Y(n3310) );
  INVX1 U437 ( .A(n3312), .Y(n422) );
  AOI22X1 U438 ( .A0(n438), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B0(n3311), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .Y(n3312) );
  AOI22X1 U439 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .A1(n418), .B0(n3317), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .Y(n3318) );
  XOR2X1 U440 ( .A(n3302), .B(n29), .Y(n3319) );
  NAND2X1 U441 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(n29) );
  AOI22X1 U442 ( .A0(n409), .A1(n412), .B0(n3301), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .Y(n3302) );
  XOR2X1 U443 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[5]) );
  XOR2X1 U444 ( .A(n418), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .Y(n3317) );
  XOR2X1 U445 ( .A(n412), .B(n409), .Y(n3301) );
  OR3XL U446 ( .A(output_previous_1[11]), .B(output_previous_1[12]), .C(n3788), 
        .Y(n3786) );
  AND2X2 U447 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer4_128126480_128126592)
         );
  AND2X2 U448 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer4_128126816_128126928)
         );
  XOR2X1 U449 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128126816_128126928)
         );
  XOR2X1 U450 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128237920_128238088)
         );
  XOR2X1 U451 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128126480_128126592)
         );
  XOR2X1 U452 ( .A(n425), .B(n3299), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128263168_128126424_128126648)
         );
  XOR2X1 U453 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .B(n3301), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128126760_128237640_128237808)
         );
  XOR2X1 U454 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .B(n3279), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128263224_128263392_128263504)
         );
  XOR2X1 U455 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .B(n3271), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128249696_128249808_128262328)
         );
  XOR2X1 U456 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .B(n3275), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128262720_128262832_128263000)
         );
  XNOR2X1 U457 ( .A(n4000), .B(n463), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[9]) );
  NOR3X1 U458 ( .A(output_previous_1[13]), .B(output_previous_1[14]), 
        .C(n3786), .Y(n3785) );
  NOR2BX1 U459 ( .AN(n3785), .B(output_previous_1[15]), .Y(n3784) );
  INVX1 U460 ( .A(output_previous_1[9]), .Y(n1210) );
  XOR2X1 U461 ( .A(n897), .B(n2829), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128262496_128126088_128126312)
         );
  XOR2X1 U462 ( .A(n1056), .B(n3063), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128262496_128126088_128126312)
         );
  XOR2X1 U463 ( .A(n579), .B(n3531), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128262496_128126088_128126312)
         );
  XOR2X1 U464 ( .A(n738), .B(n2595), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128262496_128126088_128126312)
         );
  XOR2X1 U465 ( .A(n913), .B(n906), .Y(n2827) );
  XOR2X1 U466 ( .A(n1072), .B(n1065), .Y(n3061) );
  XOR2X1 U467 ( .A(n595), .B(n588), .Y(n3529) );
  XOR2X1 U468 ( .A(n754), .B(n747), .Y(n2593) );
  XOR2X1 U469 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .B(n2827), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128125752_128125976_128126144)
         );
  XOR2X1 U470 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .B(n2593), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128125752_128125976_128126144)
         );
  BUFX3 U471 ( .A(n873), .Y(n124) );
  BUFX3 U472 ( .A(n1032), .Y(n128) );
  BUFX3 U473 ( .A(n555), .Y(n116) );
  BUFX3 U474 ( .A(n714), .Y(n120) );
  INVX1 U475 ( .A(n2828), .Y(n905) );
  AOI22X1 U476 ( .A0(n906), .A1(n913), .B0(n2827), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .Y(n2828) );
  INVX1 U477 ( .A(n3062), .Y(n1064) );
  AOI22X1 U478 ( .A0(n1065), .A1(n1072), .B0(n3061), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .Y(n3062) );
  INVX1 U479 ( .A(n3530), .Y(n587) );
  AOI22X1 U480 ( .A0(n588), .A1(n595), .B0(n3529), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .Y(n3530) );
  INVX1 U481 ( .A(n2594), .Y(n746) );
  AOI22X1 U482 ( .A0(n747), .A1(n754), .B0(n2593), 
        .B1(input_times_b0_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .Y(n2594) );
  BUFX3 U483 ( .A(n873), .Y(n123) );
  BUFX3 U484 ( .A(n1032), .Y(n127) );
  BUFX3 U485 ( .A(n555), .Y(n115) );
  BUFX3 U486 ( .A(n714), .Y(n119) );
  NOR3X1 U487 ( .A(n2311), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_8), .C(n3713), 
        .Y(n3711) );
  NOR3X1 U488 ( .A(n2332), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_8), .C(n3761), 
        .Y(n3759) );
  NOR3X1 U489 ( .A(n2374), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_8), .C(n3857), 
        .Y(n3855) );
  NOR3X1 U490 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn47), 
        .B(input_times_b0_mul_componentxunsigned_output_8), .C(n3665), 
        .Y(n3663) );
  INVX1 U491 ( .A(n2826), .Y(n914) );
  AOI22X1 U492 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .A1(n926), .B0(n2825), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .Y(n2826) );
  INVX1 U493 ( .A(n2592), .Y(n755) );
  AOI22X1 U494 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .A1(n767), .B0(n2591), 
        .B1(input_times_b0_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .Y(n2592) );
  AOI22X1 U495 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .A1(n894), .B0(n2849), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .Y(n2850) );
  INVX1 U496 ( .A(n3082), .Y(n1049) );
  AOI22X1 U497 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .A1(n1050), .B0(n3081), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .Y(n3082) );
  AOI22X1 U498 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .A1(n1053), .B0(n3083), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .Y(n3084) );
  INVX1 U499 ( .A(n3550), .Y(n572) );
  AOI22X1 U500 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .A1(n573), .B0(n3549), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .Y(n3550) );
  AOI22X1 U501 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .A1(n576), .B0(n3551), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .Y(n3552) );
  AOI22X1 U502 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .A1(n735), .B0(n2615), 
        .B1(input_times_b0_mul_componentxUMxsum_layer4_128126760_128237640_128237808), 
        .Y(n2616) );
  XOR2X1 U503 ( .A(n955), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .Y(n2819) );
  XOR2X1 U504 ( .A(n1114), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .Y(n3053) );
  XOR2X1 U505 ( .A(n637), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .Y(n3521) );
  XOR2X1 U506 ( .A(n796), 
        .B(input_times_b0_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .Y(n2585) );
  XOR2X1 U507 ( .A(n926), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .Y(n2825) );
  XOR2X1 U508 ( .A(n1085), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .Y(n3059) );
  XOR2X1 U509 ( .A(n608), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .Y(n3527) );
  XOR2X1 U510 ( .A(n767), 
        .B(input_times_b0_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .Y(n2591) );
  XOR2X1 U511 ( .A(n891), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .Y(n2847) );
  XOR2X1 U512 ( .A(n894), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .Y(n2849) );
  XOR2X1 U513 ( .A(n1050), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .Y(n3081) );
  XOR2X1 U514 ( .A(n1053), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .Y(n3083) );
  XOR2X1 U515 ( .A(n573), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .Y(n3549) );
  XOR2X1 U516 ( .A(n576), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .Y(n3551) );
  XOR2X1 U517 ( .A(n732), 
        .B(input_times_b0_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .Y(n2613) );
  XOR2X1 U518 ( .A(n735), 
        .B(input_times_b0_mul_componentxUMxcarry_layer4_128126816_128126928), 
        .Y(n2615) );
  XOR2X1 U519 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B(n941), .Y(n2837) );
  XOR2X1 U520 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B(n1100), .Y(n3071) );
  XOR2X1 U521 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B(n623), .Y(n3539) );
  XOR2X1 U522 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B(n782), .Y(n2603) );
  XOR2X1 U523 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B(n937), .Y(n2839) );
  XOR2X1 U524 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B(n1096), .Y(n3073) );
  XOR2X1 U525 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B(n619), .Y(n3541) );
  XOR2X1 U526 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B(n778), .Y(n2605) );
  XOR2X1 U527 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B(n925), .Y(n2841) );
  XOR2X1 U528 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B(n1084), .Y(n3075) );
  XOR2X1 U529 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B(n607), .Y(n3543) );
  XOR2X1 U530 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B(n766), .Y(n2607) );
  XOR2X1 U531 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B(n914), .Y(n2843) );
  XOR2X1 U532 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B(n1073), .Y(n3077) );
  XOR2X1 U533 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B(n596), .Y(n3545) );
  XOR2X1 U534 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B(n755), .Y(n2609) );
  XOR2X1 U535 ( .A(n888), .B(n885), .Y(n2833) );
  XOR2X1 U536 ( .A(n1047), .B(n1044), .Y(n3067) );
  XOR2X1 U537 ( .A(n570), .B(n567), .Y(n3535) );
  XOR2X1 U538 ( .A(n729), .B(n726), .Y(n2599) );
  AND2X2 U539 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer4_128126480_128126592)
         );
  AND2X2 U540 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer4_128126816_128126928)
         );
  AND2X2 U541 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer4_128126480_128126592)
         );
  AND2X2 U542 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer4_128126816_128126928)
         );
  AND2X2 U543 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer4_128126480_128126592)
         );
  AND2X2 U544 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer4_128126816_128126928)
         );
  AND2X2 U545 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(input_times_b0_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer4_128126480_128126592)
         );
  AND2X2 U546 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(input_times_b0_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer4_128126816_128126928)
         );
  XOR2X1 U547 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128126816_128126928)
         );
  XOR2X1 U548 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128126816_128126928)
         );
  XOR2X1 U549 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128126816_128126928)
         );
  XOR2X1 U550 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128262720_128262832_128263000), 
        .B(input_times_b0_mul_componentxUMxsum_layer3_128262216_128262384_128262552), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128126816_128126928) );
  XOR2X1 U551 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .B(n2821), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128124744_128124968_128125136)
         );
  XOR2X1 U552 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .B(n3055), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128124744_128124968_128125136)
         );
  XOR2X1 U553 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .B(n3523), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128124744_128124968_128125136)
         );
  XOR2X1 U554 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .B(n2587), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128124744_128124968_128125136)
         );
  XOR2X1 U555 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .B(n2823), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128125080_128125304_128125472)
         );
  XOR2X1 U556 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .B(n3057), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128125080_128125304_128125472)
         );
  XOR2X1 U557 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .B(n3525), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128125080_128125304_128125472)
         );
  XOR2X1 U558 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .B(n2589), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128125080_128125304_128125472)
         );
  XOR2X1 U559 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .B(n2825), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128125416_128125640_128125808)
         );
  XOR2X1 U560 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .B(n3059), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128125416_128125640_128125808)
         );
  XOR2X1 U561 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .B(n3527), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128125416_128125640_128125808)
         );
  XOR2X1 U562 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .B(n2591), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128125416_128125640_128125808)
         );
  XOR2X1 U563 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .B(n3061), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128125752_128125976_128126144)
         );
  XOR2X1 U564 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128248800_128249024_128249192), 
        .B(n3529), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128125752_128125976_128126144)
         );
  XOR2X1 U565 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128126480_128126592)
         );
  XOR2X1 U566 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128126480_128126592)
         );
  XOR2X1 U567 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128126480_128126592)
         );
  XOR2X1 U568 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128249696_128249808_128262328), 
        .B(input_times_b0_mul_componentxUMxsum_layer3_128197128_128249304_128249528), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128126480_128126592) );
  XOR2X1 U569 ( .A(n901), .B(n2831), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128263168_128126424_128126648)
         );
  XOR2X1 U570 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .B(n2833), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128126760_128237640_128237808)
         );
  XOR2X1 U571 ( .A(n1060), .B(n3065), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128263168_128126424_128126648)
         );
  XOR2X1 U572 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .B(n3067), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128126760_128237640_128237808)
         );
  XOR2X1 U573 ( .A(n583), .B(n3533), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128263168_128126424_128126648)
         );
  XOR2X1 U574 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .B(n3535), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128126760_128237640_128237808)
         );
  XOR2X1 U575 ( .A(n742), .B(n2597), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128263168_128126424_128126648)
         );
  XOR2X1 U576 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .B(n2599), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128126760_128237640_128237808)
         );
  AND2X2 U577 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219456_128219680)
         );
  AND2X2 U578 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219288_128219512)
         );
  AND2X2 U579 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219456_128219680)
         );
  AND2X2 U580 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219288_128219512)
         );
  AND2X2 U581 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219456_128219680)
         );
  AND2X2 U582 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219288_128219512)
         );
  AND2X2 U583 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(input_times_b0_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer5_128219456_128219680)
         );
  AND2X2 U584 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(input_times_b0_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer5_128219288_128219512)
         );
  AND2X2 U585 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n958), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219624_128219848)
         );
  AND2X2 U586 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n1117), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219624_128219848)
         );
  AND2X2 U587 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n640), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219624_128219848)
         );
  AND2X2 U588 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n799), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer5_128219624_128219848)
         );
  AND2X2 U589 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n949), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219792_128220016)
         );
  AND2X2 U590 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n1108), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219792_128220016)
         );
  AND2X2 U591 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n631), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219792_128220016)
         );
  AND2X2 U592 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n790), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer5_128219792_128220016)
         );
  XOR2X1 U593 ( .A(n2834), .B(n30), .Y(n2851) );
  NAND2X1 U594 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(n30) );
  AOI22X1 U595 ( .A0(n885), .A1(n888), .B0(n2833), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .Y(n2834) );
  XOR2X1 U596 ( .A(n3068), .B(n31), .Y(n3085) );
  NAND2X1 U597 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(n31) );
  AOI22X1 U598 ( .A0(n1044), .A1(n1047), .B0(n3067), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .Y(n3068) );
  XOR2X1 U599 ( .A(n3536), .B(n32), .Y(n3553) );
  NAND2X1 U600 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(n32) );
  AOI22X1 U601 ( .A0(n567), .A1(n570), .B0(n3535), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .Y(n3536) );
  XOR2X1 U602 ( .A(n2600), .B(n33), .Y(n2617) );
  NAND2X1 U603 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(input_times_b0_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(n33) );
  AOI22X1 U604 ( .A0(n726), .A1(n729), .B0(n2599), 
        .B1(input_times_b0_mul_componentxUMxsum_layer3_128262664_128262888_128263056), 
        .Y(n2600) );
  XOR2X1 U605 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128219456_128219680)
         );
  XOR2X1 U606 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128219288_128219512)
         );
  XOR2X1 U607 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128219456_128219680)
         );
  XOR2X1 U608 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128219456_128219680)
         );
  XOR2X1 U609 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128247120_128124240_128124520), 
        .B(input_times_b0_mul_componentxUMxcarry_layer4_128124072_128124296), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128219456_128219680) );
  XOR2X1 U610 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(input_times_b0_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128219288_128219512) );
  XOR2X1 U611 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .B(n2817), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128247456_128124464_128124688)
         );
  XOR2X1 U612 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .B(n2815), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128247120_128124240_128124520)
         );
  XOR2X1 U613 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .B(n3051), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128247456_128124464_128124688)
         );
  XOR2X1 U614 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .B(n3049), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128247120_128124240_128124520)
         );
  XOR2X1 U615 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .B(n3519), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128247456_128124464_128124688)
         );
  XOR2X1 U616 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .B(n3517), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128247120_128124240_128124520)
         );
  XOR2X1 U617 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .B(n2583), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128247456_128124464_128124688)
         );
  XOR2X1 U618 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .B(n2581), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128247120_128124240_128124520)
         );
  XOR2X1 U619 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128247680_128247792), 
        .B(n2819), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128124632_128124800_128124912)
         );
  XOR2X1 U620 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128247680_128247792), 
        .B(n3053), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128124632_128124800_128124912)
         );
  XOR2X1 U621 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128247680_128247792), 
        .B(n3521), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128124632_128124800_128124912)
         );
  XOR2X1 U622 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128247680_128247792), 
        .B(n2585), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128124632_128124800_128124912)
         );
  XOR2X1 U623 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n958), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128219624_128219848)
         );
  XOR2X1 U624 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n1117), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128219624_128219848)
         );
  XOR2X1 U625 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n640), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128219624_128219848)
         );
  XOR2X1 U626 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128247456_128124464_128124688), 
        .B(n799), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128219624_128219848) );
  XOR2X1 U627 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n949), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128219792_128220016)
         );
  XOR2X1 U628 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n1108), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128219792_128220016)
         );
  XOR2X1 U629 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n631), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128219792_128220016)
         );
  XOR2X1 U630 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128124632_128124800_128124912), 
        .B(n790), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128219792_128220016) );
  INVX1 U631 ( .A(n2820), .Y(n941) );
  AOI22X1 U632 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .A1(n955), .B0(n2819), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer3_128247680_128247792), 
        .Y(n2820) );
  INVX1 U633 ( .A(n3054), .Y(n1100) );
  AOI22X1 U634 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .A1(n1114), .B0(n3053), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer3_128247680_128247792), 
        .Y(n3054) );
  INVX1 U635 ( .A(n3522), .Y(n623) );
  AOI22X1 U636 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .A1(n637), .B0(n3521), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer3_128247680_128247792), 
        .Y(n3522) );
  INVX1 U637 ( .A(n2586), .Y(n782) );
  AOI22X1 U638 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer3_128222208_128247288_128247512), 
        .A1(n796), .B0(n2585), 
        .B1(input_times_b0_mul_componentxUMxsum_layer3_128247680_128247792), 
        .Y(n2586) );
  INVX1 U639 ( .A(n3060), .Y(n1073) );
  AOI22X1 U640 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .A1(n1085), .B0(n3059), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .Y(n3060) );
  INVX1 U641 ( .A(n3528), .Y(n596) );
  AOI22X1 U642 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer3_128248464_128248632), 
        .A1(n608), .B0(n3527), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer3_128248296_128248520_128248688), 
        .Y(n3528) );
  INVX1 U643 ( .A(n2848), .Y(n890) );
  AOI22X1 U644 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .A1(n891), .B0(n2847), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .Y(n2848) );
  INVX1 U645 ( .A(n2614), .Y(n731) );
  AOI22X1 U646 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer4_128126480_128126592), 
        .A1(n732), .B0(n2613), 
        .B1(input_times_b0_mul_componentxUMxsum_layer4_128263168_128126424_128126648), 
        .Y(n2614) );
  INVX1 U647 ( .A(n2838), .Y(n929) );
  AOI22X1 U648 ( .A0(n941), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B0(n2837), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .Y(n2838) );
  INVX1 U649 ( .A(n3072), .Y(n1088) );
  AOI22X1 U650 ( .A0(n1100), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B0(n3071), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .Y(n3072) );
  INVX1 U651 ( .A(n3540), .Y(n611) );
  AOI22X1 U652 ( .A0(n623), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B0(n3539), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .Y(n3540) );
  INVX1 U653 ( .A(n2604), .Y(n770) );
  AOI22X1 U654 ( .A0(n782), 
        .A1(input_times_b0_mul_componentxUMxsum_layer3_128248016_128248128), 
        .B0(n2603), 
        .B1(input_times_b0_mul_componentxUMxsum_layer4_128124744_128124968_128125136), 
        .Y(n2604) );
  INVX1 U655 ( .A(n2840), .Y(n916) );
  AOI22X1 U656 ( .A0(n937), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B0(n2839), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .Y(n2840) );
  INVX1 U657 ( .A(n3074), .Y(n1075) );
  AOI22X1 U658 ( .A0(n1096), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B0(n3073), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .Y(n3074) );
  INVX1 U659 ( .A(n3542), .Y(n598) );
  AOI22X1 U660 ( .A0(n619), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B0(n3541), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .Y(n3542) );
  INVX1 U661 ( .A(n2606), .Y(n757) );
  AOI22X1 U662 ( .A0(n778), 
        .A1(input_times_b0_mul_componentxUMxsum_layer3_128248464_128248632), 
        .B0(n2605), 
        .B1(input_times_b0_mul_componentxUMxsum_layer4_128125080_128125304_128125472), 
        .Y(n2606) );
  INVX1 U663 ( .A(n2842), .Y(n907) );
  AOI22X1 U664 ( .A0(n925), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B0(n2841), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .Y(n2842) );
  INVX1 U665 ( .A(n3076), .Y(n1066) );
  AOI22X1 U666 ( .A0(n1084), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B0(n3075), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .Y(n3076) );
  INVX1 U667 ( .A(n3544), .Y(n589) );
  AOI22X1 U668 ( .A0(n607), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B0(n3543), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .Y(n3544) );
  INVX1 U669 ( .A(n2608), .Y(n748) );
  AOI22X1 U670 ( .A0(n766), 
        .A1(input_times_b0_mul_componentxUMxsum_layer3_128248856_128248968_128249136), 
        .B0(n2607), 
        .B1(input_times_b0_mul_componentxUMxsum_layer4_128125416_128125640_128125808), 
        .Y(n2608) );
  INVX1 U671 ( .A(n2844), .Y(n898) );
  AOI22X1 U672 ( .A0(n914), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B0(n2843), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .Y(n2844) );
  INVX1 U673 ( .A(n3078), .Y(n1057) );
  AOI22X1 U674 ( .A0(n1073), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B0(n3077), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .Y(n3078) );
  INVX1 U675 ( .A(n3546), .Y(n580) );
  AOI22X1 U676 ( .A0(n596), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B0(n3545), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .Y(n3546) );
  INVX1 U677 ( .A(n2610), .Y(n739) );
  AOI22X1 U678 ( .A0(n755), 
        .A1(input_times_b0_mul_componentxUMxsum_layer3_128249360_128249472_128249640), 
        .B0(n2609), 
        .B1(input_times_b0_mul_componentxUMxsum_layer4_128125752_128125976_128126144), 
        .Y(n2610) );
  XOR2X1 U679 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[5]) );
  XOR2X1 U680 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[5]) );
  XOR2X1 U681 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[5]) );
  XOR2X1 U682 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(input_times_b0_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[5]) );
  XOR2X1 U683 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128237920_128238088)
         );
  XOR2X1 U684 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128237920_128238088)
         );
  XOR2X1 U685 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128237920_128238088)
         );
  XOR2X1 U686 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128263672_128263840), 
        .B(input_times_b0_mul_componentxUMxsum_layer3_128263224_128263392_128263504), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128237920_128238088) );
  AND2X2 U687 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer5_128219120_128219344)
         );
  AND2X2 U688 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer5_128219120_128219344)
         );
  AND2X2 U689 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer5_128219120_128219344)
         );
  AND2X2 U690 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128123904_128124128), 
        .B(input_times_b0_mul_componentxUMxcarry_layer4_128123792_128123960), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer5_128219120_128219344)
         );
  XOR2X1 U691 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128219288_128219512)
         );
  XOR2X1 U692 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128124072_128124296), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer4_128123904_128124128), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128219288_128219512)
         );
  XNOR2X1 U693 ( .A(n3914), .B(n940), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[9]) );
  XNOR2X1 U694 ( .A(n3957), .B(n1099), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[9]) );
  XNOR2X1 U695 ( .A(n4043), .B(n622), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[9]) );
  XNOR2X1 U696 ( .A(n3871), .B(n781), 
        .Y(input_times_b0_div_componentxinput_A_inverted[9]) );
  NAND3X1 U697 ( .A(output_previous_1[11]), .B(output_previous_1[10]), 
        .C(output_previous_1[12]), .Y(output_contracterxn5) );
  OR3XL U698 ( .A(output_previous_1[12]), .B(output_previous_1[13]), 
        .C(output_previous_1[14]), .Y(output_contracterxn8) );
  INVX1 U699 ( .A(n3250), .Y(n489) );
  AOI22X1 U700 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .A1(n497), .B0(n3249), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_127827304_127827416), 
        .Y(n3250) );
  XOR2X1 U701 ( .A(n497), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .Y(n3249) );
  XOR2X1 U702 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B(n489), .Y(n3283) );
  XOR2X1 U703 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B(n482), .Y(n3285) );
  INVX1 U704 ( .A(n232), .Y(n398) );
  BUFX3 U705 ( .A(n1203), .Y(n134) );
  INVX1 U706 ( .A(n3284), .Y(n481) );
  AOI22X1 U707 ( .A0(n489), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B0(n3283), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .Y(n3284) );
  BUFX3 U708 ( .A(n1203), .Y(n133) );
  NOR3X1 U709 ( .A(n480), .B(n473), .C(n4001), .Y(n4000) );
  NOR3X1 U710 ( .A(n423), .B(n417), .C(n4008), .Y(n4007) );
  INVX1 U711 ( .A(n3254), .Y(n478) );
  AOI22X1 U712 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .A1(n483), .B0(n3253), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .Y(n3254) );
  INVX1 U713 ( .A(n3260), .Y(n449) );
  AOI22X1 U714 ( .A0(n451), .A1(n457), .B0(n3259), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .Y(n3260) );
  INVX1 U715 ( .A(n3262), .Y(n437) );
  AOI22X1 U716 ( .A0(n439), .A1(n447), .B0(n3261), 
        .B1(output_p1_times_a1_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .Y(n3262) );
  NAND3BX1 U717 ( .AN(n453), .B(n4547), .C(n4000), .Y(n4009) );
  NOR2BX1 U718 ( .AN(n4007), .B(n408), .Y(n4006) );
  OR3XL U719 ( .A(\output_signal[3] ), .B(\output_signal[4] ), .C(n3781), 
        .Y(n3779) );
  XOR2X1 U720 ( .A(n471), .B(n3255), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128222208_128247288_128247512)
         );
  XOR2X1 U721 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .B(n3215), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128223440_128223608_128223776)
         );
  XOR2X1 U722 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .B(n3221), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128224280_128224448_128224560)
         );
  XOR2X1 U723 ( .A(n483), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .Y(n3253) );
  XOR2X1 U724 ( .A(n470), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .Y(n3289) );
  XOR2X1 U725 ( .A(n459), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .Y(n3291) );
  XOR2X1 U726 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .Y(n3263) );
  XOR2X1 U727 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .Y(n3267) );
  XOR2X1 U728 ( .A(n457), .B(n451), .Y(n3259) );
  XOR2X1 U729 ( .A(n447), .B(n439), .Y(n3261) );
  XOR2X1 U730 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B(n433), .Y(n3297) );
  OR3XL U731 ( .A(n441), .B(n432), .C(n4009), .Y(n4008) );
  OR3XL U732 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[5]), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[6]), .C(n3811), 
        .Y(n3809) );
  AND2X2 U733 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer3_128247680_128247792)
         );
  AND2X2 U734 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer3_128248016_128248128)
         );
  AND2X2 U735 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer3_128248464_128248632)
         );
  XOR2X1 U736 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128248016_128248128)
         );
  XOR2X1 U737 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .B(n3263), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128248856_128248968_128249136)
         );
  XOR2X1 U738 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .B(n3251), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128246616_128246840_128247008)
         );
  XOR2X1 U739 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .B(n3253), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128246952_128247176_128247344)
         );
  XOR2X1 U740 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128247680_128247792)
         );
  XOR2X1 U741 ( .A(n461), .B(n3257), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128222880_128247624_128247848)
         );
  XOR2X1 U742 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .B(n3259), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128247960_128248184_128248352)
         );
  XOR2X1 U743 ( 
        .A(output_p1_times_a1_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .B(n3261), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128248296_128248520_128248688)
         );
  XOR2X1 U744 ( .A(n456), .B(n3265), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128248800_128249024_128249192)
         );
  AND2X2 U745 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer3_128246000_128246168)
         );
  AND2X2 U746 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer4_128123904_128124128)
         );
  AND2X2 U747 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer4_128123792_128123960)
         );
  AND2X2 U748 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n496), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer4_128124072_128124296)
         );
  NAND2BX1 U749 ( .AN(n401), .B(n4006), .Y(n4005) );
  XOR2X1 U750 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128123904_128124128)
         );
  XOR2X1 U751 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127827304_127827416), 
        .B(n3249), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128246504_128246672_128246784)
         );
  XOR2X1 U752 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .B(n3247), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_127827080_128246280_128246560)
         );
  XOR2X1 U753 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n496), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128124072_128124296)
         );
  INVX1 U754 ( .A(n3290), .Y(n460) );
  AOI22X1 U755 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .A1(n470), .B0(n3289), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .Y(n3290) );
  INVX1 U756 ( .A(n3292), .Y(n448) );
  AOI22X1 U757 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .A1(n459), .B0(n3291), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .Y(n3292) );
  INVX1 U758 ( .A(n3264), .Y(n430) );
  AOI22X1 U759 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B0(n3263), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .Y(n3264) );
  XNOR2X1 U760 ( .A(n4007), .B(n408), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[15]) );
  XNOR2X1 U761 ( .A(n4006), .B(n401), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[16]) );
  XOR2X1 U762 ( .A(n4008), .B(n423), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[13]) );
  XNOR2X1 U763 ( .A(n34), .B(n417), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[14]) );
  NOR2X1 U764 ( .A(n423), .B(n4008), .Y(n34) );
  INVX1 U765 ( .A(n3298), .Y(n415) );
  AOI22X1 U766 ( .A0(n433), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B0(n3297), .B1(n421), .Y(n3298) );
  INVX1 U767 ( .A(n3268), .Y(n421) );
  AOI22X1 U768 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B0(n3267), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .Y(n3268) );
  INVX1 U769 ( .A(n3286), .Y(n472) );
  AOI22X1 U770 ( .A0(n482), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B0(n3285), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .Y(n3286) );
  INVX1 U771 ( .A(n3300), .Y(n418) );
  AOI22X1 U772 ( .A0(n419), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B0(n3299), .B1(n425), .Y(n3300) );
  XOR2X1 U773 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[3]) );
  XOR2X1 U774 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[4]) );
  XOR2X1 U775 ( .A(n454), .B(n3237), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128197464_128197688_128197856)
         );
  XOR2X1 U776 ( .A(n475), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .Y(n3271) );
  XOR2X1 U777 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .Y(n3235) );
  XOR2X1 U778 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .Y(n3275) );
  XOR2X1 U779 ( 
        .A(output_p1_times_a1_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .Y(n3279) );
  XOR2X1 U780 ( .A(n428), .B(n455), .Y(n3219) );
  XOR2X1 U781 ( .A(n426), .B(n446), .Y(n3225) );
  XOR2X1 U782 ( .A(n444), .B(n403), .Y(n3237) );
  XOR2X1 U783 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B(n419), .Y(n3299) );
  XOR2X1 U784 ( .A(n424), .B(n442), .Y(n3273) );
  OR3XL U785 ( .A(n495), .B(n488), .C(n4002), .Y(n4001) );
  XOR2X1 U786 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128248464_128248632)
         );
  XOR2X1 U787 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .B(n3267), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128249360_128249472_128249640)
         );
  XOR2X1 U788 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .B(n3227), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128224952_128225120_128225232)
         );
  XOR2X1 U789 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .B(n3235), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128197520_128197632_128197800)
         );
  XOR2X1 U790 ( .A(n406), .B(n3277), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128262664_128262888_128263056)
         );
  OR3XL U791 ( .A(n509), .B(n503), .C(n4003), .Y(n4002) );
  XOR2X1 U792 ( .A(n420), .B(n3269), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128197128_128249304_128249528)
         );
  XOR2X1 U793 ( .A(n413), .B(n3273), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128262216_128262384_128262552)
         );
  INVX1 U794 ( .A(n4547), .Y(n463) );
  XOR2X1 U795 ( .A(n3238), .B(n3240), .Y(n3281) );
  AOI22X1 U796 ( .A0(n403), .A1(n444), .B0(n3237), .B1(n454), .Y(n3238) );
  INVX1 U797 ( .A(n3276), .Y(n409) );
  AOI22X1 U798 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B0(n3275), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .Y(n3276) );
  XOR2X1 U799 ( .A(n4009), .B(n441), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[11]) );
  XNOR2X1 U800 ( .A(n35), .B(n432), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[12]) );
  NOR2X1 U801 ( .A(n4009), .B(n441), .Y(n35) );
  XOR2X1 U802 ( .A(n4010), .B(n453), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[10]) );
  NAND2X1 U803 ( .A(n4000), .B(n4547), .Y(n4010) );
  INVX1 U804 ( .A(n3274), .Y(n412) );
  AOI22X1 U805 ( .A0(n442), .A1(n424), .B0(n3273), .B1(n413), .Y(n3274) );
  INVX1 U806 ( .A(n3272), .Y(n425) );
  AOI22X1 U807 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .A1(n475), .B0(n3271), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .Y(n3272) );
  XOR2X1 U808 ( .A(n4177), .B(n4178), .Y(output_previous_1[13]) );
  XOR2X1 U809 ( .A(n4181), .B(n4182), .Y(output_previous_1[11]) );
  XOR2X1 U810 ( .A(n4176), .B(n4175), .Y(output_previous_1[14]) );
  XOR2X1 U811 ( .A(n4154), .B(n4155), .Y(output_previous_1[8]) );
  XOR2X1 U812 ( .A(n4184), .B(n4183), .Y(output_previous_1[10]) );
  XOR2X1 U813 ( .A(n4180), .B(n4179), .Y(output_previous_1[12]) );
  XOR2X1 U814 ( .A(n4152), .B(n4153), .Y(output_previous_1[9]) );
  AOI22X1 U815 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .A1(output_p1_times_a1_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B0(n3279), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .Y(n3280) );
  XOR2X1 U816 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .Y(n3241) );
  XOR2X1 U817 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .B(n3239), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128198080_128198192_128198360)
         );
  XOR2X1 U818 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128263672_128263840)
         );
  XOR2X1 U819 ( .A(n4001), .B(n480), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[7]) );
  XNOR2X1 U820 ( .A(n36), .B(n473), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[8]) );
  NOR2X1 U821 ( .A(n480), .B(n4001), .Y(n36) );
  XOR2X1 U822 ( 
        .A(output_p1_times_a1_mul_componentxUMxcarry_layer3_128263672_128263840), 
        .B(n3303), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128237752_128237976_128238144)
         );
  AND2X2 U823 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer3_128263672_128263840)
         );
  XOR2X1 U824 ( .A(n404), .B(n402), .Y(n3303) );
  INVX1 U825 ( .A(n3280), .Y(n402) );
  INVX1 U826 ( .A(n3236), .Y(n406) );
  AOI22X1 U827 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B0(n3235), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .Y(n3236) );
  XOR2X1 U828 ( .A(n4173), .B(n4174), .Y(output_previous_1[15]) );
  XOR2X1 U829 ( .A(n4171), .B(n1205), .Y(output_previous_1[16]) );
  XOR2X1 U830 ( .A(n4002), .B(n495), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[5]) );
  XNOR2X1 U831 ( .A(n37), .B(n503), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[4]) );
  NOR2X1 U832 ( .A(n509), .B(n4003), .Y(n37) );
  XNOR2X1 U833 ( .A(n38), .B(n488), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[6]) );
  NOR2X1 U834 ( .A(n495), .B(n4002), .Y(n38) );
  BUFX3 U835 ( .A(n80), .Y(n114) );
  BUFX3 U836 ( .A(n80), .Y(n113) );
  XOR2X1 U837 ( .A(n4003), .B(n509), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[3]) );
  INVX1 U838 ( .A(n2796), .Y(n906) );
  AOI22X1 U839 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B0(n2795), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .Y(n2796) );
  INVX1 U840 ( .A(n2562), .Y(n747) );
  AOI22X1 U841 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .A1(input_times_b0_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B0(n2561), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .Y(n2562) );
  XOR2X1 U842 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .Y(n2795) );
  XOR2X1 U843 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .Y(n3029) );
  XOR2X1 U844 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .Y(n3497) );
  XOR2X1 U845 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .Y(n2561) );
  XOR2X1 U846 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B(n909), .Y(n2829) );
  XOR2X1 U847 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B(n1068), .Y(n3063) );
  XOR2X1 U848 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B(n591), .Y(n3531) );
  XOR2X1 U849 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B(n750), .Y(n2595) );
  INVX1 U850 ( .A(n190), .Y(n873) );
  INVX1 U851 ( .A(n211), .Y(n1032) );
  INVX1 U852 ( .A(n253), .Y(n555) );
  INVX1 U853 ( .A(n281), .Y(n714) );
  INVX1 U854 ( .A(n3030), .Y(n1065) );
  AOI22X1 U855 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B0(n3029), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .Y(n3030) );
  INVX1 U856 ( .A(n3498), .Y(n588) );
  AOI22X1 U857 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer2_128223440_128223608_128223776), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer2_127715424_128223048_128223272), 
        .B0(n3497), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .Y(n3498) );
  NOR3X1 U858 ( .A(n899), .B(n893), .C(n3922), .Y(n3921) );
  NOR3X1 U859 ( .A(n1058), .B(n1052), .C(n3965), .Y(n3964) );
  NOR3X1 U860 ( .A(n581), .B(n575), .C(n4051), .Y(n4050) );
  NOR3X1 U861 ( .A(n740), .B(n734), .C(n3879), .Y(n3878) );
  INVX1 U862 ( .A(n2786), .Y(n955) );
  AOI22X1 U863 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .A1(n960), .B0(n2785), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .Y(n2786) );
  INVX1 U864 ( .A(n3020), .Y(n1114) );
  AOI22X1 U865 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .A1(n1119), .B0(n3019), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .Y(n3020) );
  INVX1 U866 ( .A(n3488), .Y(n637) );
  AOI22X1 U867 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .A1(n642), .B0(n3487), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .Y(n3488) );
  INVX1 U868 ( .A(n2552), .Y(n796) );
  AOI22X1 U869 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .A1(n801), .B0(n2551), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .Y(n2552) );
  INVX1 U870 ( .A(n2822), .Y(n937) );
  AOI22X1 U871 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .A1(n947), .B0(n2821), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .Y(n2822) );
  INVX1 U872 ( .A(n2588), .Y(n778) );
  AOI22X1 U873 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .A1(n788), .B0(n2587), 
        .B1(input_times_b0_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .Y(n2588) );
  INVX1 U874 ( .A(n2824), .Y(n925) );
  AOI22X1 U875 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .A1(n936), .B0(n2823), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .Y(n2824) );
  INVX1 U876 ( .A(n2794), .Y(n913) );
  AOI22X1 U877 ( .A0(n915), .A1(n924), .B0(n2793), 
        .B1(input_p1_times_b1_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .Y(n2794) );
  INVX1 U878 ( .A(n2590), .Y(n766) );
  AOI22X1 U879 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .A1(n777), .B0(n2589), 
        .B1(input_times_b0_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .Y(n2590) );
  INVX1 U880 ( .A(n2560), .Y(n754) );
  AOI22X1 U881 ( .A0(n756), .A1(n765), .B0(n2559), 
        .B1(input_times_b0_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .Y(n2560) );
  INVX1 U882 ( .A(n2808), .Y(n885) );
  AOI22X1 U883 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B0(n2807), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .Y(n2808) );
  INVX1 U884 ( .A(n2574), .Y(n726) );
  AOI22X1 U885 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .A1(input_times_b0_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B0(n2573), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .Y(n2574) );
  INVX1 U886 ( .A(n2830), .Y(n891) );
  AOI22X1 U887 ( .A0(n909), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B0(n2829), .B1(n897), .Y(n2830) );
  INVX1 U888 ( .A(n2832), .Y(n894) );
  AOI22X1 U889 ( .A0(n895), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B0(n2831), .B1(n901), .Y(n2832) );
  INVX1 U890 ( .A(n3040), .Y(n1047) );
  AOI22X1 U891 ( .A0(n1077), .A1(n1059), .B0(n3039), .B1(n1048), .Y(n3040) );
  INVX1 U892 ( .A(n3508), .Y(n570) );
  AOI22X1 U893 ( .A0(n600), .A1(n582), .B0(n3507), .B1(n571), .Y(n3508) );
  INVX1 U894 ( .A(n2596), .Y(n732) );
  AOI22X1 U895 ( .A0(n750), 
        .A1(input_times_b0_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B0(n2595), .B1(n738), .Y(n2596) );
  INVX1 U896 ( .A(n2598), .Y(n735) );
  AOI22X1 U897 ( .A0(n736), 
        .A1(input_times_b0_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B0(n2597), .B1(n742), .Y(n2598) );
  NAND3BX1 U898 ( .AN(n930), .B(n4441), .C(n3914), .Y(n3923) );
  NAND3BX1 U899 ( .AN(n1089), .B(n4494), .C(n3957), .Y(n3966) );
  NAND3BX1 U900 ( .AN(n612), .B(n4600), .C(n4043), .Y(n4052) );
  NAND3BX1 U901 ( .AN(n771), .B(input_times_b0_mul_componentxn90), .C(n3871), 
        .Y(n3880) );
  NOR2BX1 U902 ( .AN(n3921), .B(n884), .Y(n3920) );
  NOR2BX1 U903 ( .AN(n3964), .B(n1043), .Y(n3963) );
  NOR2BX1 U904 ( .AN(n4050), .B(n566), .Y(n4049) );
  NOR2BX1 U905 ( .AN(n3878), .B(n725), .Y(n3877) );
  XOR2X1 U906 ( .A(n948), .B(n2787), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128222208_128247288_128247512)
         );
  XOR2X1 U907 ( .A(n1107), .B(n3021), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128222208_128247288_128247512)
         );
  XOR2X1 U908 ( .A(n630), .B(n3489), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128222208_128247288_128247512)
         );
  XOR2X1 U909 ( .A(n789), .B(n2553), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128222208_128247288_128247512)
         );
  XOR2X1 U910 ( .A(n974), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .Y(n2781) );
  XOR2X1 U911 ( .A(n1133), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .Y(n3015) );
  XOR2X1 U912 ( .A(n656), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .Y(n3483) );
  XOR2X1 U913 ( .A(n815), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .Y(n2547) );
  XOR2X1 U914 ( .A(n960), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .Y(n2785) );
  XOR2X1 U915 ( .A(n1119), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .Y(n3019) );
  XOR2X1 U916 ( .A(n642), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .Y(n3487) );
  XOR2X1 U917 ( .A(n801), 
        .B(input_times_b0_mul_componentxUMxcarry_layer2_127827752_127827920), 
        .Y(n2551) );
  XOR2X1 U918 ( .A(n947), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .Y(n2821) );
  XOR2X1 U919 ( .A(n936), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .Y(n2823) );
  XOR2X1 U920 ( .A(n1106), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .Y(n3055) );
  XOR2X1 U921 ( .A(n1095), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .Y(n3057) );
  XOR2X1 U922 ( .A(n629), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .Y(n3523) );
  XOR2X1 U923 ( .A(n618), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .Y(n3525) );
  XOR2X1 U924 ( .A(n788), 
        .B(input_times_b0_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .Y(n2587) );
  XOR2X1 U925 ( .A(n777), 
        .B(input_times_b0_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .Y(n2589) );
  XOR2X1 U926 ( .A(n952), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .Y(n2803) );
  XOR2X1 U927 ( .A(n1111), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .Y(n3037) );
  XOR2X1 U928 ( .A(n634), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .Y(n3505) );
  XOR2X1 U929 ( .A(n793), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .Y(n2569) );
  XOR2X1 U930 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .Y(n2799) );
  XOR2X1 U931 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .Y(n3033) );
  XOR2X1 U932 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .Y(n3501) );
  XOR2X1 U933 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .Y(n2565) );
  XOR2X1 U934 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .Y(n2807) );
  XOR2X1 U935 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .Y(n3041) );
  XOR2X1 U936 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .Y(n3509) );
  XOR2X1 U937 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .Y(n2573) );
  XOR2X1 U938 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B(n966), .Y(n2815) );
  XOR2X1 U939 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B(n1125), .Y(n3049) );
  XOR2X1 U940 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B(n648), .Y(n3517) );
  XOR2X1 U941 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B(n807), .Y(n2581) );
  XOR2X1 U942 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B(n959), .Y(n2817) );
  XOR2X1 U943 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B(n1118), .Y(n3051) );
  XOR2X1 U944 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B(n641), .Y(n3519) );
  XOR2X1 U945 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B(n800), .Y(n2583) );
  XOR2X1 U946 ( .A(n934), .B(n928), .Y(n2791) );
  XOR2X1 U947 ( .A(n1093), .B(n1087), .Y(n3025) );
  XOR2X1 U948 ( .A(n616), .B(n610), .Y(n3493) );
  XOR2X1 U949 ( .A(n775), .B(n769), .Y(n2557) );
  XOR2X1 U950 ( .A(n924), .B(n915), .Y(n2793) );
  XOR2X1 U951 ( .A(n1083), .B(n1074), .Y(n3027) );
  XOR2X1 U952 ( .A(n606), .B(n597), .Y(n3495) );
  XOR2X1 U953 ( .A(n765), .B(n756), .Y(n2559) );
  XOR2X1 U954 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B(n895), .Y(n2831) );
  XOR2X1 U955 ( .A(n900), .B(n918), .Y(n2805) );
  XOR2X1 U956 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B(n1054), .Y(n3065) );
  XOR2X1 U957 ( .A(n1059), .B(n1077), .Y(n3039) );
  XOR2X1 U958 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B(n577), .Y(n3533) );
  XOR2X1 U959 ( .A(n582), .B(n600), .Y(n3507) );
  XOR2X1 U960 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B(n736), .Y(n2597) );
  XOR2X1 U961 ( .A(n741), .B(n759), .Y(n2571) );
  OR3XL U962 ( .A(n917), .B(n908), .C(n3923), .Y(n3922) );
  OR3XL U963 ( .A(n1076), .B(n1067), .C(n3966), .Y(n3965) );
  OR3XL U964 ( .A(n599), .B(n590), .C(n4052), .Y(n4051) );
  OR3XL U965 ( .A(n758), .B(n749), .C(n3880), .Y(n3879) );
  AND2X2 U966 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer3_128248016_128248128)
         );
  AND2X2 U967 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer3_128247680_128247792)
         );
  AND2X2 U968 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer3_128248016_128248128)
         );
  AND2X2 U969 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer3_128247680_128247792)
         );
  AND2X2 U970 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer3_128248016_128248128)
         );
  AND2X2 U971 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer3_128247680_128247792)
         );
  AND2X2 U972 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer3_128248016_128248128)
         );
  AND2X2 U973 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer3_128247680_128247792)
         );
  AND2X2 U974 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer3_128248464_128248632)
         );
  AND2X2 U975 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer3_128248464_128248632)
         );
  AND2X2 U976 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer3_128248464_128248632)
         );
  AND2X2 U977 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer3_128248464_128248632)
         );
  XOR2X1 U978 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128248464_128248632)
         );
  XOR2X1 U979 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128248464_128248632)
         );
  XOR2X1 U980 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128248464_128248632)
         );
  XOR2X1 U981 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128223384_128223552), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128222936_128223104_128223216), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128248464_128248632) );
  XOR2X1 U982 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .B(n2795), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128248856_128248968_128249136)
         );
  XOR2X1 U983 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .B(n3029), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128248856_128248968_128249136)
         );
  XOR2X1 U984 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .B(n3497), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128248856_128248968_128249136)
         );
  XOR2X1 U985 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128223888_128224112_128224056), 
        .B(n2561), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128248856_128248968_128249136)
         );
  XOR2X1 U986 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .B(n2799), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128249360_128249472_128249640)
         );
  XOR2X1 U987 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .B(n3033), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128249360_128249472_128249640)
         );
  XOR2X1 U988 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .B(n3501), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128249360_128249472_128249640)
         );
  XOR2X1 U989 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .B(n2565), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128249360_128249472_128249640)
         );
  XOR2X1 U990 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .B(n2783), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128246616_128246840_128247008)
         );
  XOR2X1 U991 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .B(n3017), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128246616_128246840_128247008)
         );
  XOR2X1 U992 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .B(n3485), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128246616_128246840_128247008)
         );
  XOR2X1 U993 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .B(n2549), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128246616_128246840_128247008)
         );
  XOR2X1 U994 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .B(n2785), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128246952_128247176_128247344)
         );
  XOR2X1 U995 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .B(n3019), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128246952_128247176_128247344)
         );
  XOR2X1 U996 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .B(n3487), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128246952_128247176_128247344)
         );
  XOR2X1 U997 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127827584_127827808_128221256), 
        .B(n2551), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128246952_128247176_128247344)
         );
  XOR2X1 U998 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128247680_128247792)
         );
  XOR2X1 U999 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128247680_128247792)
         );
  XOR2X1 U1000 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128247680_128247792)
         );
  XOR2X1 U1001 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128221760_128221928_128222040), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_127635584_128221368_128221592), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128247680_128247792) );
  XOR2X1 U1002 ( .A(n938), .B(n2789), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128222880_128247624_128247848)
         );
  XOR2X1 U1003 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .B(n2791), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128247960_128248184_128248352)
         );
  XOR2X1 U1004 ( .A(n1097), .B(n3023), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128222880_128247624_128247848)
         );
  XOR2X1 U1005 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .B(n3025), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128247960_128248184_128248352)
         );
  XOR2X1 U1006 ( .A(n620), .B(n3491), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128222880_128247624_128247848)
         );
  XOR2X1 U1007 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .B(n3493), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128247960_128248184_128248352)
         );
  XOR2X1 U1008 ( .A(n779), .B(n2555), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128222880_128247624_128247848)
         );
  XOR2X1 U1009 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .B(n2557), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128247960_128248184_128248352)
         );
  XOR2X1 U1010 ( 
        .A(input_p1_times_b1_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .B(n2793), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128248296_128248520_128248688)
         );
  XOR2X1 U1011 ( 
        .A(input_p2_times_b2_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .B(n3027), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128248296_128248520_128248688)
         );
  XOR2X1 U1012 ( 
        .A(output_p2_times_a2_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .B(n3495), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128248296_128248520_128248688)
         );
  XOR2X1 U1013 ( 
        .A(input_times_b0_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .B(n2559), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128248296_128248520_128248688)
         );
  XOR2X1 U1014 ( .A(n933), .B(n2797), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128248800_128249024_128249192)
         );
  XOR2X1 U1015 ( .A(n1092), .B(n3031), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128248800_128249024_128249192)
         );
  XOR2X1 U1016 ( .A(n615), .B(n3499), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128248800_128249024_128249192)
         );
  XOR2X1 U1017 ( .A(n774), .B(n2563), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128248800_128249024_128249192)
         );
  XOR2X1 U1018 ( .A(n896), .B(n2801), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128197128_128249304_128249528)
         );
  XOR2X1 U1019 ( .A(n889), .B(n2805), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128262216_128262384_128262552)
         );
  XOR2X1 U1020 ( .A(n1055), .B(n3035), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128197128_128249304_128249528)
         );
  XOR2X1 U1021 ( .A(n1048), .B(n3039), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128262216_128262384_128262552)
         );
  XOR2X1 U1022 ( .A(n578), .B(n3503), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128197128_128249304_128249528)
         );
  XOR2X1 U1023 ( .A(n571), .B(n3507), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128262216_128262384_128262552)
         );
  XOR2X1 U1024 ( .A(n737), .B(n2567), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128197128_128249304_128249528)
         );
  XOR2X1 U1025 ( .A(n730), .B(n2571), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128262216_128262384_128262552)
         );
  AND2X2 U1026 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer4_128123904_128124128)
         );
  AND2X2 U1027 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer4_128123904_128124128)
         );
  AND2X2 U1028 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer4_128123904_128124128)
         );
  AND2X2 U1029 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(input_times_b0_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer4_128123904_128124128)
         );
  AND2X2 U1030 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n973), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer4_128124072_128124296)
         );
  AND2X2 U1031 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n1132), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer4_128124072_128124296)
         );
  AND2X2 U1032 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n655), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer4_128124072_128124296)
         );
  AND2X2 U1033 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n814), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer4_128124072_128124296)
         );
  NAND2BX1 U1034 ( .AN(n876), .B(n3920), .Y(n3919) );
  NAND2BX1 U1035 ( .AN(n1035), .B(n3963), .Y(n3962) );
  NAND2BX1 U1036 ( .AN(n558), .B(n4049), .Y(n4048) );
  NAND2BX1 U1037 ( .AN(n717), .B(n3877), .Y(n3876) );
  XOR2X1 U1038 ( .A(n875), 
        .B(input_p1_times_b1_mul_componentxUMxsecond_vector[17]), .Y(n2313) );
  XOR2X1 U1039 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer5_128315744_128315968_128316136), 
        .B(n2856), .Y(input_p1_times_b1_mul_componentxUMxsecond_vector[17]) );
  INVX1 U1040 ( .A(n2855), .Y(n875) );
  XOR2X1 U1041 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128237752_128237976_128238144), 
        .B(n2851), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer5_128315744_128315968_128316136)
         );
  XOR2X1 U1042 ( .A(n1034), 
        .B(input_p2_times_b2_mul_componentxUMxsecond_vector[17]), .Y(n2334) );
  XOR2X1 U1043 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer5_128315744_128315968_128316136), 
        .B(n3090), .Y(input_p2_times_b2_mul_componentxUMxsecond_vector[17]) );
  INVX1 U1044 ( .A(n3089), .Y(n1034) );
  XOR2X1 U1045 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128237752_128237976_128238144), 
        .B(n3085), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer5_128315744_128315968_128316136)
         );
  XOR2X1 U1046 ( .A(n557), 
        .B(output_p2_times_a2_mul_componentxUMxsecond_vector[17]), .Y(n2376)
         );
  XOR2X1 U1047 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer5_128315744_128315968_128316136), 
        .B(n3558), .Y(output_p2_times_a2_mul_componentxUMxsecond_vector[17])
         );
  INVX1 U1048 ( .A(n3557), .Y(n557) );
  XOR2X1 U1049 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128237752_128237976_128238144), 
        .B(n3553), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer5_128315744_128315968_128316136)
         );
  XOR2X1 U1050 ( .A(n716), 
        .B(input_times_b0_mul_componentxUMxsecond_vector[17]), 
        .Y(input_times_b0_mul_componentxUMxAdder_finalxn475) );
  XOR2X1 U1051 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer5_128315744_128315968_128316136), 
        .B(n2622), .Y(input_times_b0_mul_componentxUMxsecond_vector[17]) );
  INVX1 U1052 ( .A(n2621), .Y(n716) );
  XOR2X1 U1053 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128237752_128237976_128238144), 
        .B(n2617), 
        .Y(input_times_b0_mul_componentxUMxsum_layer5_128315744_128315968_128316136)
         );
  XOR2X1 U1054 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127827304_127827416), 
        .B(n2781), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128246504_128246672_128246784)
         );
  XOR2X1 U1055 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .B(n2779), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_127827080_128246280_128246560)
         );
  XOR2X1 U1056 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127827304_127827416), 
        .B(n3015), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128246504_128246672_128246784)
         );
  XOR2X1 U1057 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .B(n3013), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_127827080_128246280_128246560)
         );
  XOR2X1 U1058 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127827304_127827416), 
        .B(n3483), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128246504_128246672_128246784)
         );
  XOR2X1 U1059 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .B(n3481), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_127827080_128246280_128246560)
         );
  XOR2X1 U1060 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127827304_127827416), 
        .B(n2547), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128246504_128246672_128246784)
         );
  XOR2X1 U1061 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .B(n2545), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_127827080_128246280_128246560)
         );
  XOR2X1 U1062 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .B(n2803), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128249696_128249808_128262328)
         );
  XOR2X1 U1063 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .B(n2807), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128262720_128262832_128263000)
         );
  XOR2X1 U1064 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .B(n3037), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128249696_128249808_128262328)
         );
  XOR2X1 U1065 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .B(n3041), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128262720_128262832_128263000)
         );
  XOR2X1 U1066 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .B(n3505), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128249696_128249808_128262328)
         );
  XOR2X1 U1067 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .B(n3509), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128262720_128262832_128263000)
         );
  XOR2X1 U1068 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .B(n2569), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128249696_128249808_128262328)
         );
  XOR2X1 U1069 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .B(n2573), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128262720_128262832_128263000)
         );
  XOR2X1 U1070 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n973), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128124072_128124296)
         );
  XOR2X1 U1071 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n1132), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128124072_128124296)
         );
  XOR2X1 U1072 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n655), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128124072_128124296)
         );
  XOR2X1 U1073 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128246504_128246672_128246784), 
        .B(n814), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128124072_128124296) );
  INVX1 U1074 ( .A(n2782), .Y(n966) );
  AOI22X1 U1075 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .A1(n974), .B0(n2781), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_127827304_127827416), 
        .Y(n2782) );
  INVX1 U1076 ( .A(n3016), .Y(n1125) );
  AOI22X1 U1077 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .A1(n1133), .B0(n3015), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_127827304_127827416), 
        .Y(n3016) );
  INVX1 U1078 ( .A(n3484), .Y(n648) );
  AOI22X1 U1079 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .A1(n656), .B0(n3483), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_127827304_127827416), 
        .Y(n3484) );
  INVX1 U1080 ( .A(n2548), .Y(n807) );
  AOI22X1 U1081 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer2_127731808_127826912_127827136), 
        .A1(n815), .B0(n2547), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_127827304_127827416), 
        .Y(n2548) );
  INVX1 U1082 ( .A(n3056), .Y(n1096) );
  AOI22X1 U1083 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .A1(n1106), .B0(n3055), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .Y(n3056) );
  INVX1 U1084 ( .A(n3524), .Y(n619) );
  AOI22X1 U1085 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer3_128247680_128247792), 
        .A1(n629), .B0(n3523), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer3_128222880_128247624_128247848), 
        .Y(n3524) );
  INVX1 U1086 ( .A(n3058), .Y(n1084) );
  AOI22X1 U1087 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .A1(n1095), .B0(n3057), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .Y(n3058) );
  INVX1 U1088 ( .A(n3526), .Y(n607) );
  AOI22X1 U1089 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer3_128248016_128248128), 
        .A1(n618), .B0(n3525), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer3_128247960_128248184_128248352), 
        .Y(n3526) );
  INVX1 U1090 ( .A(n3042), .Y(n1044) );
  AOI22X1 U1091 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B0(n3041), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .Y(n3042) );
  INVX1 U1092 ( .A(n3510), .Y(n567) );
  AOI22X1 U1093 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer2_128197016_128197240_128197352), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer2_127627392_128196680_128196848), 
        .B0(n3509), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_128197520_128197632_128197800), 
        .Y(n3510) );
  XNOR2X1 U1094 ( .A(n3921), .B(n884), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[15]) );
  XNOR2X1 U1095 ( .A(n3964), .B(n1043), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[15]) );
  XNOR2X1 U1096 ( .A(n4050), .B(n566), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[15]) );
  XNOR2X1 U1097 ( .A(n3878), .B(n725), 
        .Y(input_times_b0_div_componentxinput_A_inverted[15]) );
  XNOR2X1 U1098 ( .A(n3920), .B(n876), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[16]) );
  XNOR2X1 U1099 ( .A(n3963), .B(n1035), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[16]) );
  XNOR2X1 U1100 ( .A(n4049), .B(n558), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[16]) );
  XNOR2X1 U1101 ( .A(n3877), .B(n717), 
        .Y(input_times_b0_div_componentxinput_A_inverted[16]) );
  XNOR2X1 U1102 ( .A(n39), .B(n893), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[14]) );
  NOR2X1 U1103 ( .A(n899), .B(n3922), .Y(n39) );
  XNOR2X1 U1104 ( .A(n40), .B(n1052), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[14]) );
  NOR2X1 U1105 ( .A(n1058), .B(n3965), .Y(n40) );
  XNOR2X1 U1106 ( .A(n41), .B(n575), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[14]) );
  NOR2X1 U1107 ( .A(n581), .B(n4051), .Y(n41) );
  XNOR2X1 U1108 ( .A(n42), .B(n734), 
        .Y(input_times_b0_div_componentxinput_A_inverted[14]) );
  NOR2X1 U1109 ( .A(n740), .B(n3879), .Y(n42) );
  INVX1 U1110 ( .A(n2792), .Y(n926) );
  AOI22X1 U1111 ( .A0(n928), .A1(n934), .B0(n2791), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .Y(n2792) );
  INVX1 U1112 ( .A(n3026), .Y(n1085) );
  AOI22X1 U1113 ( .A0(n1087), .A1(n1093), .B0(n3025), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .Y(n3026) );
  INVX1 U1114 ( .A(n3494), .Y(n608) );
  AOI22X1 U1115 ( .A0(n610), .A1(n616), .B0(n3493), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .Y(n3494) );
  INVX1 U1116 ( .A(n2558), .Y(n767) );
  AOI22X1 U1117 ( .A0(n769), .A1(n775), .B0(n2557), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_128222376_128222600_128222768), 
        .Y(n2558) );
  INVX1 U1118 ( .A(n3028), .Y(n1072) );
  AOI22X1 U1119 ( .A0(n1074), .A1(n1083), .B0(n3027), 
        .B1(input_p2_times_b2_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .Y(n3028) );
  INVX1 U1120 ( .A(n3496), .Y(n595) );
  AOI22X1 U1121 ( .A0(n597), .A1(n606), .B0(n3495), 
        .B1(output_p2_times_a2_mul_componentxUMxcarry_layer2_128223384_128223552), 
        .Y(n3496) );
  INVX1 U1122 ( .A(n2806), .Y(n888) );
  AOI22X1 U1123 ( .A0(n918), .A1(n900), .B0(n2805), .B1(n889), .Y(n2806) );
  INVX1 U1124 ( .A(n3064), .Y(n1050) );
  AOI22X1 U1125 ( .A0(n1068), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B0(n3063), .B1(n1056), .Y(n3064) );
  INVX1 U1126 ( .A(n3066), .Y(n1053) );
  AOI22X1 U1127 ( .A0(n1054), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B0(n3065), .B1(n1060), .Y(n3066) );
  INVX1 U1128 ( .A(n3532), .Y(n573) );
  AOI22X1 U1129 ( .A0(n591), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer2_128196792_128196960_128197184), 
        .B0(n3531), .B1(n579), .Y(n3532) );
  INVX1 U1130 ( .A(n3534), .Y(n576) );
  AOI22X1 U1131 ( .A0(n577), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer2_128198024_128197968), 
        .B0(n3533), .B1(n583), .Y(n3534) );
  INVX1 U1132 ( .A(n2572), .Y(n729) );
  AOI22X1 U1133 ( .A0(n759), .A1(n741), .B0(n2571), .B1(n730), .Y(n2572) );
  INVX1 U1134 ( .A(n2800), .Y(n897) );
  AOI22X1 U1135 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B0(n2799), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .Y(n2800) );
  INVX1 U1136 ( .A(n2804), .Y(n901) );
  AOI22X1 U1137 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .A1(n952), .B0(n2803), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .Y(n2804) );
  INVX1 U1138 ( .A(n3034), .Y(n1056) );
  AOI22X1 U1139 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B0(n3033), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .Y(n3034) );
  INVX1 U1140 ( .A(n3038), .Y(n1060) );
  AOI22X1 U1141 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .A1(n1111), .B0(n3037), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .Y(n3038) );
  INVX1 U1142 ( .A(n3502), .Y(n579) );
  AOI22X1 U1143 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B0(n3501), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .Y(n3502) );
  INVX1 U1144 ( .A(n3506), .Y(n583) );
  AOI22X1 U1145 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .A1(n634), .B0(n3505), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .Y(n3506) );
  INVX1 U1146 ( .A(n2566), .Y(n738) );
  AOI22X1 U1147 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer2_128224280_128224448_128224560), 
        .A1(input_times_b0_mul_componentxUMxsum_layer2_128223720_128223944_128224168), 
        .B0(n2565), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_128224728_128224896_128225064), 
        .Y(n2566) );
  INVX1 U1148 ( .A(n2570), .Y(n742) );
  AOI22X1 U1149 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer2_128224392_128224616_128224784), 
        .A1(n793), .B0(n2569), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_128224952_128225120_128225232), 
        .Y(n2570) );
  INVX1 U1150 ( .A(n2816), .Y(n958) );
  AOI22X1 U1151 ( .A0(n966), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B0(n2815), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .Y(n2816) );
  INVX1 U1152 ( .A(n3050), .Y(n1117) );
  AOI22X1 U1153 ( .A0(n1125), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B0(n3049), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .Y(n3050) );
  INVX1 U1154 ( .A(n3518), .Y(n640) );
  AOI22X1 U1155 ( .A0(n648), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B0(n3517), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .Y(n3518) );
  INVX1 U1156 ( .A(n2582), .Y(n799) );
  AOI22X1 U1157 ( .A0(n807), 
        .A1(input_times_b0_mul_componentxUMxsum_layer2_127827752_127827920), 
        .B0(n2581), 
        .B1(input_times_b0_mul_componentxUMxsum_layer3_128246616_128246840_128247008), 
        .Y(n2582) );
  INVX1 U1158 ( .A(n2818), .Y(n949) );
  AOI22X1 U1159 ( .A0(n959), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B0(n2817), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .Y(n2818) );
  INVX1 U1160 ( .A(n3052), .Y(n1108) );
  AOI22X1 U1161 ( .A0(n1118), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B0(n3051), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .Y(n3052) );
  INVX1 U1162 ( .A(n3520), .Y(n631) );
  AOI22X1 U1163 ( .A0(n641), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B0(n3519), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .Y(n3520) );
  INVX1 U1164 ( .A(n2584), .Y(n790) );
  AOI22X1 U1165 ( .A0(n800), 
        .A1(input_times_b0_mul_componentxUMxsum_layer2_128221424_128221536_128221704), 
        .B0(n2583), 
        .B1(input_times_b0_mul_componentxUMxsum_layer3_128246952_128247176_128247344), 
        .Y(n2584) );
  NOR3X1 U1166 ( .A(n957), .B(n950), .C(n3915), .Y(n3914) );
  NOR3X1 U1167 ( .A(n1116), .B(n1109), .C(n3958), .Y(n3957) );
  NOR3X1 U1168 ( .A(n639), .B(n632), .C(n4044), .Y(n4043) );
  NOR3X1 U1169 ( .A(n798), .B(n791), .C(n3872), .Y(n3871) );
  XOR2X1 U1170 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[4]) );
  XOR2X1 U1171 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[4]) );
  XOR2X1 U1172 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[4]) );
  XOR2X1 U1173 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(input_times_b0_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[4]) );
  XOR2X1 U1174 ( 
        .A(input_p1_times_b1_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .Y(n2811) );
  XOR2X1 U1175 ( 
        .A(input_p2_times_b2_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .Y(n3045) );
  XOR2X1 U1176 ( 
        .A(output_p2_times_a2_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .Y(n3513) );
  XOR2X1 U1177 ( 
        .A(input_times_b0_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .Y(n2577) );
  OR3XL U1178 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[5]), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[6]), .C(n3715), 
        .Y(n3713) );
  OR3XL U1179 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[5]), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[6]), .C(n3763), 
        .Y(n3761) );
  OR3XL U1180 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[5]), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[6]), .C(n3859), 
        .Y(n3857) );
  OR3XL U1181 ( .A(input_times_b0_mul_componentxUMxfirst_vector[5]), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[6]), .C(n3667), 
        .Y(n3665) );
  OR3XL U1182 ( .A(n972), .B(n965), .C(n3916), .Y(n3915) );
  OR3XL U1183 ( .A(n1131), .B(n1124), .C(n3959), .Y(n3958) );
  OR3XL U1184 ( .A(n654), .B(n647), .C(n4045), .Y(n4044) );
  OR3XL U1185 ( .A(n813), .B(n806), .C(n3873), .Y(n3872) );
  XOR2X1 U1186 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128248016_128248128)
         );
  XOR2X1 U1187 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128248016_128248128)
         );
  XOR2X1 U1188 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128248016_128248128)
         );
  XOR2X1 U1189 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128222432_128222544_128222712), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128221872_128222096_128222264), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128248016_128248128) );
  XOR2X1 U1190 ( .A(n882), .B(n2809), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128262664_128262888_128263056)
         );
  XOR2X1 U1191 ( .A(n1041), .B(n3043), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128262664_128262888_128263056)
         );
  XOR2X1 U1192 ( .A(n564), .B(n3511), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128262664_128262888_128263056)
         );
  XOR2X1 U1193 ( .A(n723), .B(n2575), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128262664_128262888_128263056)
         );
  XOR2X1 U1194 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .B(n2811), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128263224_128263392_128263504)
         );
  XOR2X1 U1195 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .B(n3045), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128263224_128263392_128263504)
         );
  XOR2X1 U1196 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .B(n3513), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128263224_128263392_128263504)
         );
  XOR2X1 U1197 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .B(n2577), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128263224_128263392_128263504)
         );
  AND2X2 U1198 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer3_128246000_128246168)
         );
  AND2X2 U1199 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer3_128246000_128246168)
         );
  AND2X2 U1200 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer3_128246000_128246168)
         );
  AND2X2 U1201 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(input_times_b0_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer3_128246000_128246168)
         );
  AND2X2 U1202 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer4_128123792_128123960)
         );
  AND2X2 U1203 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer4_128123792_128123960)
         );
  AND2X2 U1204 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer4_128123792_128123960)
         );
  AND2X2 U1205 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128246112_128246336), 
        .B(input_times_b0_mul_componentxUMxcarry_layer3_128246000_128246168), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer4_128123792_128123960)
         );
  XOR2X1 U1206 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128123904_128124128)
         );
  XOR2X1 U1207 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128123904_128124128)
         );
  XOR2X1 U1208 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128123904_128124128)
         );
  XOR2X1 U1209 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_127827080_128246280_128246560), 
        .B(input_times_b0_mul_componentxUMxcarry_layer3_128246112_128246336), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128123904_128124128) );
  XOR2X1 U1210 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128263672_128263840)
         );
  XOR2X1 U1211 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128263672_128263840)
         );
  XOR2X1 U1212 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128263672_128263840)
         );
  XOR2X1 U1213 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128263672_128263840) );
  XOR2X1 U1214 ( .A(n3923), .B(n917), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[11]) );
  XOR2X1 U1215 ( .A(n3966), .B(n1076), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[11]) );
  XOR2X1 U1216 ( .A(n4052), .B(n599), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[11]) );
  XOR2X1 U1217 ( .A(n3880), .B(n758), 
        .Y(input_times_b0_div_componentxinput_A_inverted[11]) );
  XOR2X1 U1218 ( .A(n3922), .B(n899), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[13]) );
  XOR2X1 U1219 ( .A(n3965), .B(n1058), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[13]) );
  XOR2X1 U1220 ( .A(n4051), .B(n581), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[13]) );
  XOR2X1 U1221 ( .A(n3879), .B(n740), 
        .Y(input_times_b0_div_componentxinput_A_inverted[13]) );
  XNOR2X1 U1222 ( .A(n43), .B(n908), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[12]) );
  NOR2X1 U1223 ( .A(n3923), .B(n917), .Y(n43) );
  XNOR2X1 U1224 ( .A(n44), .B(n1067), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[12]) );
  NOR2X1 U1225 ( .A(n3966), .B(n1076), .Y(n44) );
  XNOR2X1 U1226 ( .A(n45), .B(n590), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[12]) );
  NOR2X1 U1227 ( .A(n4052), .B(n599), .Y(n45) );
  XNOR2X1 U1228 ( .A(n46), .B(n749), 
        .Y(input_times_b0_div_componentxinput_A_inverted[12]) );
  NOR2X1 U1229 ( .A(n3880), .B(n758), .Y(n46) );
  XOR2X1 U1230 ( .A(n3924), .B(n930), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[10]) );
  NAND2X1 U1231 ( .A(n3914), .B(n4441), .Y(n3924) );
  XOR2X1 U1232 ( .A(n3967), .B(n1089), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[10]) );
  NAND2X1 U1233 ( .A(n3957), .B(n4494), .Y(n3967) );
  XOR2X1 U1234 ( .A(n4053), .B(n612), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[10]) );
  NAND2X1 U1235 ( .A(n4043), .B(n4600), .Y(n4053) );
  XOR2X1 U1236 ( .A(n3881), .B(n771), 
        .Y(input_times_b0_div_componentxinput_A_inverted[10]) );
  NAND2X1 U1237 ( .A(n3871), .B(input_times_b0_mul_componentxn90), .Y(n3881)
         );
  XOR2X1 U1238 ( 
        .A(input_p1_times_b1_mul_componentxUMxcarry_layer3_128263672_128263840), 
        .B(n2835), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128237752_128237976_128238144)
         );
  AND2X2 U1239 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer3_128263672_128263840)
         );
  XOR2X1 U1240 ( .A(n880), .B(n878), .Y(n2835) );
  INVX1 U1241 ( .A(n2810), .Y(n880) );
  XOR2X1 U1242 ( 
        .A(input_p2_times_b2_mul_componentxUMxcarry_layer3_128263672_128263840), 
        .B(n3069), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128237752_128237976_128238144)
         );
  AND2X2 U1243 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer3_128263672_128263840)
         );
  XOR2X1 U1244 ( .A(n1039), .B(n1037), .Y(n3069) );
  INVX1 U1245 ( .A(n3044), .Y(n1039) );
  XOR2X1 U1246 ( 
        .A(output_p2_times_a2_mul_componentxUMxcarry_layer3_128263672_128263840), 
        .B(n3537), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128237752_128237976_128238144)
         );
  AND2X2 U1247 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer3_128263672_128263840)
         );
  XOR2X1 U1248 ( .A(n562), .B(n560), .Y(n3537) );
  INVX1 U1249 ( .A(n3512), .Y(n562) );
  XOR2X1 U1250 ( 
        .A(input_times_b0_mul_componentxUMxcarry_layer3_128263672_128263840), 
        .B(n2601), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128237752_128237976_128238144)
         );
  AND2X2 U1251 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128198976_128199144), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128198472_128198640_128198808), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer3_128263672_128263840)
         );
  XOR2X1 U1252 ( .A(n721), .B(n719), .Y(n2601) );
  INVX1 U1253 ( .A(n2576), .Y(n721) );
  INVX1 U1254 ( .A(n2812), .Y(n878) );
  AOI22X1 U1255 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .A1(input_p1_times_b1_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B0(n2811), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .Y(n2812) );
  INVX1 U1256 ( .A(n3046), .Y(n1037) );
  AOI22X1 U1257 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .A1(input_p2_times_b2_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B0(n3045), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .Y(n3046) );
  INVX1 U1258 ( .A(n3514), .Y(n560) );
  AOI22X1 U1259 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .A1(output_p2_times_a2_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B0(n3513), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .Y(n3514) );
  INVX1 U1260 ( .A(n2578), .Y(n719) );
  AOI22X1 U1261 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer2_128197464_128197688_128197856), 
        .A1(input_times_b0_mul_componentxUMxcarry_layer2_128198024_128197968), 
        .B0(n2577), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_128198080_128198192_128198360), 
        .Y(n2578) );
  XOR2X1 U1262 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[3]) );
  XOR2X1 U1263 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[3]) );
  XOR2X1 U1264 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[3]) );
  XOR2X1 U1265 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127672448_127826240_127826520), 
        .B(input_times_b0_mul_componentxUMxcarry_layer2_127826128_127826296), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[3]) );
  OR3XL U1266 ( .A(n986), .B(n980), .C(n3917), .Y(n3916) );
  OR3XL U1267 ( .A(n1145), .B(n1139), .C(n3960), .Y(n3959) );
  OR3XL U1268 ( .A(n668), .B(n662), .C(n4046), .Y(n4045) );
  OR3XL U1269 ( .A(n827), .B(n821), .C(n3874), .Y(n3873) );
  INVX1 U1270 ( .A(n4441), .Y(n940) );
  INVX1 U1271 ( .A(n4494), .Y(n1099) );
  INVX1 U1272 ( .A(n4600), .Y(n622) );
  INVX1 U1273 ( .A(input_times_b0_mul_componentxn90), .Y(n781) );
  XOR2X1 U1274 ( .A(n3915), .B(n957), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[7]) );
  XOR2X1 U1275 ( .A(n3958), .B(n1116), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[7]) );
  XOR2X1 U1276 ( .A(n4044), .B(n639), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[7]) );
  XOR2X1 U1277 ( .A(n3872), .B(n798), 
        .Y(input_times_b0_div_componentxinput_A_inverted[7]) );
  XNOR2X1 U1278 ( .A(n47), .B(n950), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[8]) );
  NOR2X1 U1279 ( .A(n957), .B(n3915), .Y(n47) );
  XNOR2X1 U1280 ( .A(n48), .B(n1109), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[8]) );
  NOR2X1 U1281 ( .A(n1116), .B(n3958), .Y(n48) );
  XNOR2X1 U1282 ( .A(n49), .B(n632), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[8]) );
  NOR2X1 U1283 ( .A(n639), .B(n4044), .Y(n49) );
  XNOR2X1 U1284 ( .A(n50), .B(n791), 
        .Y(input_times_b0_div_componentxinput_A_inverted[8]) );
  NOR2X1 U1285 ( .A(n798), .B(n3872), .Y(n50) );
  XOR2X1 U1286 ( .A(n3916), .B(n972), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[5]) );
  XOR2X1 U1287 ( .A(n3959), .B(n1131), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[5]) );
  XOR2X1 U1288 ( .A(n4045), .B(n654), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[5]) );
  XOR2X1 U1289 ( .A(n3873), .B(n813), 
        .Y(input_times_b0_div_componentxinput_A_inverted[5]) );
  XNOR2X1 U1290 ( .A(n51), .B(n965), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[6]) );
  NOR2X1 U1291 ( .A(n972), .B(n3916), .Y(n51) );
  XNOR2X1 U1292 ( .A(n52), .B(n1124), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[6]) );
  NOR2X1 U1293 ( .A(n1131), .B(n3959), .Y(n52) );
  XNOR2X1 U1294 ( .A(n53), .B(n647), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[6]) );
  NOR2X1 U1295 ( .A(n654), .B(n4045), .Y(n53) );
  XNOR2X1 U1296 ( .A(n54), .B(n806), 
        .Y(input_times_b0_div_componentxinput_A_inverted[6]) );
  NOR2X1 U1297 ( .A(n813), .B(n3873), .Y(n54) );
  BUFX3 U1298 ( .A(n81), .Y(n126) );
  BUFX3 U1299 ( .A(n82), .Y(n130) );
  BUFX3 U1300 ( .A(n83), .Y(n118) );
  BUFX3 U1301 ( .A(n84), .Y(n122) );
  BUFX3 U1302 ( .A(n81), .Y(n125) );
  BUFX3 U1303 ( .A(n82), .Y(n129) );
  BUFX3 U1304 ( .A(n83), .Y(n117) );
  BUFX3 U1305 ( .A(n84), .Y(n121) );
  XOR2X1 U1306 ( .A(n3917), .B(n986), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[3]) );
  XOR2X1 U1307 ( .A(n3960), .B(n1145), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[3]) );
  XOR2X1 U1308 ( .A(n4046), .B(n668), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[3]) );
  XOR2X1 U1309 ( .A(n3874), .B(n827), 
        .Y(input_times_b0_div_componentxinput_A_inverted[3]) );
  XNOR2X1 U1310 ( .A(n55), .B(n980), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[4]) );
  NOR2X1 U1311 ( .A(n986), .B(n3917), .Y(n55) );
  XNOR2X1 U1312 ( .A(n56), .B(n1139), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[4]) );
  NOR2X1 U1313 ( .A(n1145), .B(n3960), .Y(n56) );
  XNOR2X1 U1314 ( .A(n57), .B(n662), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[4]) );
  NOR2X1 U1315 ( .A(n668), .B(n4046), .Y(n57) );
  XNOR2X1 U1316 ( .A(n58), .B(n821), 
        .Y(input_times_b0_div_componentxinput_A_inverted[4]) );
  NOR2X1 U1317 ( .A(n827), .B(n3874), .Y(n58) );
  NAND3BX1 U1318 ( .AN(output_contracterxn6), .B(output_previous_1[8]), 
        .C(output_previous_1[9]), .Y(output_contracterxn3) );
  NAND3BX1 U1319 ( .AN(output_contracterxn5), .B(output_previous_1[13]), 
        .C(output_previous_1[14]), .Y(output_contracterxn4) );
  NOR3X1 U1320 ( .A(output_contracterxn8), .B(output_previous_1[11]), 
        .C(output_previous_1[10]), .Y(output_contracterxn1) );
  NOR3X1 U1321 ( .A(results_a1_a2[7]), .B(results_a1_a2[8]), 
        .C(results_a1_a2_inv_inverterxn4), .Y(results_a1_a2_inv_inverterxn2)
         );
  AOI22X1 U1322 ( .A0(results_a1_a2_inv[3]), .A1(results_b0_b1_b2[3]), 
        .B0(n4164), .B1(n4165), .Y(n4163) );
  AOI22X1 U1323 ( .A0(results_a1_a2_inv[5]), .A1(results_b0_b1_b2[5]), 
        .B0(n4160), .B1(n4161), .Y(n4159) );
  AOI22X1 U1324 ( .A0(results_a1_a2_inv[7]), .A1(results_b0_b1_b2[7]), 
        .B0(n4156), .B1(n4157), .Y(n4155) );
  AOI22X1 U1325 ( .A0(results_a1_a2_inv[9]), .A1(results_b0_b1_b2[9]), 
        .B0(n4152), .B1(n4153), .Y(n4183) );
  AOI22X1 U1326 ( .A0(results_a1_a2_inv[11]), .A1(results_b0_b1_b2[11]), 
        .B0(n4181), .B1(n4182), .Y(n4179) );
  AOI22X1 U1327 ( .A0(results_a1_a2_inv[13]), .A1(results_b0_b1_b2[13]), 
        .B0(n4177), .B1(n4178), .Y(n4175) );
  OAI2BB2X1 U1328 ( .B0(n4167), .B1(n4166), .A0N(results_a1_a2_inv[2]), 
        .A1N(results_b0_b1_b2[2]), .Y(n4164) );
  OAI2BB2X1 U1329 ( .B0(n4163), .B1(n4162), .A0N(results_a1_a2_inv[4]), 
        .A1N(results_b0_b1_b2[4]), .Y(n4160) );
  OAI2BB2X1 U1330 ( .B0(n4159), .B1(n4158), .A0N(results_a1_a2_inv[6]), 
        .A1N(results_b0_b1_b2[6]), .Y(n4156) );
  OAI2BB2X1 U1331 ( .B0(n4155), .B1(n4154), .A0N(results_a1_a2_inv[8]), 
        .A1N(results_b0_b1_b2[8]), .Y(n4152) );
  OAI2BB2X1 U1332 ( .B0(n4183), .B1(n4184), .A0N(results_a1_a2_inv[10]), 
        .A1N(results_b0_b1_b2[10]), .Y(n4181) );
  OAI2BB2X1 U1333 ( .B0(n4179), .B1(n4180), .A0N(results_a1_a2_inv[12]), 
        .A1N(results_b0_b1_b2[12]), .Y(n4177) );
  OAI2BB2X1 U1334 ( .B0(n4175), .B1(n4176), .A0N(results_a1_a2_inv[14]), 
        .A1N(results_b0_b1_b2[14]), .Y(n4173) );
  INVX1 U1335 ( .A(n3192), .Y(n497) );
  AOI22X1 U1336 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .A1(n501), .B0(n3191), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .Y(n3192) );
  XNOR2X1 U1337 ( .A(results_a1_a2_inv_inverterxn2), .B(results_a1_a2[9]), 
        .Y(results_a1_a2_inv[9]) );
  XOR2X1 U1338 ( .A(n513), .B(n3193), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127731808_127826912_127827136)
         );
  XOR2X1 U1339 ( .A(results_b0_b1_b2[3]), .B(results_a1_a2_inv[3]), .Y(n4165)
         );
  XOR2X1 U1340 ( .A(results_b0_b1_b2[5]), .B(results_a1_a2_inv[5]), .Y(n4161)
         );
  XOR2X1 U1341 ( .A(results_b0_b1_b2[7]), .B(results_a1_a2_inv[7]), .Y(n4157)
         );
  XOR2X1 U1342 ( .A(results_b0_b1_b2[9]), .B(results_a1_a2_inv[9]), .Y(n4153)
         );
  XOR2X1 U1343 ( .A(results_b0_b1_b2[11]), .B(results_a1_a2_inv[11]), 
        .Y(n4182) );
  XOR2X1 U1344 ( .A(results_b0_b1_b2[13]), .B(results_a1_a2_inv[13]), 
        .Y(n4178) );
  XOR2X1 U1345 ( .A(results_b0_b1_b2[15]), .B(results_a1_a2_inv[15]), 
        .Y(n4174) );
  XOR2X1 U1346 ( .A(n501), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .Y(n3191) );
  XOR2X1 U1347 ( .A(n493), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .Y(n3251) );
  OR3XL U1348 ( .A(results_a1_a2[5]), .B(results_a1_a2[6]), 
        .C(results_a1_a2_inv_inverterxn6), .Y(results_a1_a2_inv_inverterxn4)
         );
  BUFX3 U1349 ( .A(n4557), .Y(n232) );
  AOI22X1 U1350 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_17), 
        .A1(n113), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[17]), 
        .B1(n4548), .Y(n4557) );
  XOR2X1 U1351 ( .A(n3815), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_17), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[17]) );
  XOR2X1 U1352 ( .A(n2354), .B(n2355), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_17) );
  XNOR2X1 U1353 ( .A(results_b0_b1_b2[2]), .B(results_a1_a2_inv[2]), .Y(n4166)
         );
  XNOR2X1 U1354 ( .A(results_b0_b1_b2[4]), .B(results_a1_a2_inv[4]), .Y(n4162)
         );
  XNOR2X1 U1355 ( .A(results_b0_b1_b2[6]), .B(results_a1_a2_inv[6]), .Y(n4158)
         );
  XNOR2X1 U1356 ( .A(results_b0_b1_b2[8]), .B(results_a1_a2_inv[8]), .Y(n4154)
         );
  XNOR2X1 U1357 ( .A(results_b0_b1_b2[10]), .B(results_a1_a2_inv[10]), 
        .Y(n4184) );
  XNOR2X1 U1358 ( .A(results_b0_b1_b2[12]), .B(results_a1_a2_inv[12]), 
        .Y(n4180) );
  XNOR2X1 U1359 ( .A(results_b0_b1_b2[14]), .B(results_a1_a2_inv[14]), 
        .Y(n4176) );
  BUFX3 U1360 ( .A(n4546), .Y(n231) );
  AOI22X1 U1361 ( .A0(\output_signal[0] ), .A1(n133), .B0(\output_signal[0] ), 
        .B1(n165), .Y(n4546) );
  BUFX3 U1362 ( .A(n4538), .Y(n230) );
  AOI22XL U1363 ( .A0(\output_signal[1] ), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_1_), .B1(n165), 
        .Y(n4538) );
  XOR2X1 U1364 ( .A(\output_signal[1] ), .B(\output_signal[0] ), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_1_) );
  INVX1 U1365 ( .A(n165), .Y(n1203) );
  INVX1 U1366 ( .A(n4172), .Y(n1205) );
  AOI22X1 U1367 ( .A0(results_a1_a2_inv[15]), .A1(results_b0_b1_b2[15]), 
        .B0(n4173), .B1(n4174), .Y(n4172) );
  INVX1 U1368 ( .A(n3252), .Y(n482) );
  AOI22X1 U1369 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .A1(n493), .B0(n3251), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .Y(n3252) );
  AOI22X1 U1370 ( .A0(output_previous_1[10]), .A1(n133), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_10_), .B1(n165), 
        .Y(n4545) );
  XOR2X1 U1371 ( .A(n3790), .B(output_previous_1[10]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_10_) );
  NAND2X1 U1372 ( .A(n3775), .B(n1210), .Y(n3790) );
  AOI22X1 U1373 ( .A0(output_previous_1[11]), .A1(n133), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_11_), .B1(n165), 
        .Y(n4544) );
  XOR2X1 U1374 ( .A(n3788), .B(output_previous_1[11]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_11_) );
  AOI22X1 U1375 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_9), 
        .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[9]), 
        .B1(n4548), .Y(n4547) );
  XNOR2X1 U1376 ( .A(n3807), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_9), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[9]) );
  NOR3X1 U1377 ( .A(results_a1_a2[13]), .B(results_a1_a2[14]), 
        .C(results_a1_a2_inv_inverterxn13), .Y(results_a1_a2_inv_inverterxn12)
         );
  INVX1 U1378 ( .A(n3122), .Y(n450) );
  AOI22X1 U1379 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b9), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b10), .B0(n3121), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b8), .Y(n3122) );
  INVX1 U1380 ( .A(n4561), .Y(n423) );
  AOI22X1 U1381 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_13), 
        .A1(n113), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[13]), 
        .B1(n4548), .Y(n4561) );
  XOR2X1 U1382 ( .A(n3818), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_13), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[13]) );
  INVX1 U1383 ( .A(n4558), .Y(n401) );
  AOI22X1 U1384 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_16), 
        .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[16]), 
        .B1(n4548), .Y(n4558) );
  XNOR2X1 U1385 ( .A(n3816), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_16), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[16]) );
  INVX1 U1386 ( .A(n3204), .Y(n461) );
  AOI22X1 U1387 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .A1(n512), .B0(n3203), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .Y(n3204) );
  INVX1 U1388 ( .A(n3216), .Y(n434) );
  AOI22X1 U1389 ( .A0(n511), .A1(n491), .B0(n3215), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .Y(n3216) );
  INVX1 U1390 ( .A(n3218), .Y(n456) );
  AOI22X1 U1391 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B0(n3217), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .Y(n3218) );
  INVX1 U1392 ( .A(n3116), .Y(n458) );
  AOI22X1 U1393 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b8), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b9), .B0(n3115), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b7), .Y(n3116) );
  INVX1 U1394 ( .A(n3206), .Y(n457) );
  AOI22X1 U1395 ( .A0(n486), .A1(n458), .B0(n3205), .B1(n505), .Y(n3206) );
  NAND3BX1 U1396 ( .AN(results_a1_a2[10]), .B(n1302), 
        .C(results_a1_a2_inv_inverterxn2), .Y(results_a1_a2_inv_inverterxn15)
         );
  NOR2BX1 U1397 ( .AN(results_a1_a2_inv_inverterxn12), .B(results_a1_a2[15]), 
        .Y(results_a1_a2_inv_inverterxn11) );
  XNOR2X1 U1398 ( .A(results_a1_a2_inv_inverterxn12), .B(results_a1_a2[15]), 
        .Y(results_a1_a2_inv[15]) );
  XNOR2X1 U1399 ( .A(results_a1_a2_inv_inverterxn11), .B(results_a1_a2[16]), 
        .Y(results_a1_a2_inv[16]) );
  XOR2X1 U1400 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b11), .B(n3143), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831568_127845824_127847728)
         );
  XOR2X1 U1401 ( .A(results_a1_a2_inv_inverterxn15), .B(results_a1_a2[11]), 
        .Y(results_a1_a2_inv[11]) );
  XOR2X1 U1402 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b7), .B(n3115), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831120_127845376_127847280)
         );
  XOR2X1 U1403 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b9), .B(n3127), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831344_127845600_127847504)
         );
  XOR2X1 U1404 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b10), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b9), .Y(n3121) );
  XOR2X1 U1405 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b11), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b10), .Y(n3127) );
  XOR2X1 U1406 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b12), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b11), .Y(n3135) );
  XOR2X1 U1407 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b13), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b12), .Y(n3143) );
  XOR2X1 U1408 ( .A(results_a1_a2_inv_inverterxn13), .B(results_a1_a2[13]), 
        .Y(results_a1_a2_inv[13]) );
  XOR2X1 U1409 ( .A(results_a1_a2_inv_inverterxn4), .B(results_a1_a2[7]), 
        .Y(results_a1_a2_inv[7]) );
  XOR2X1 U1410 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b8), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b7), .Y(n3109) );
  XOR2X1 U1411 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b9), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b8), .Y(n3115) );
  XOR2X1 U1412 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b9), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b8), .Y(n3137) );
  XOR2X1 U1413 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b8), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b7), .Y(n3129) );
  XOR2X1 U1414 ( .A(results_a1_a2_inv_inverterxn8), .B(results_a1_a2[3]), 
        .Y(results_a1_a2_inv[3]) );
  XOR2X1 U1415 ( .A(results_a1_a2_inv_inverterxn6), .B(results_a1_a2[5]), 
        .Y(results_a1_a2_inv[5]) );
  XOR2X1 U1416 ( .A(n508), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .Y(n3189) );
  XOR2X1 U1417 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .Y(n3199) );
  XOR2X1 U1418 ( .A(n512), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .Y(n3203) );
  XOR2X1 U1419 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .Y(n3207) );
  XOR2X1 U1420 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .Y(n3217) );
  XOR2X1 U1421 ( .A(n504), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .Y(n3221) );
  XOR2X1 U1422 ( 
        .A(output_p1_times_a1_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .Y(n3211) );
  XOR2X1 U1423 ( .A(n479), .B(n500), .Y(n3197) );
  XOR2X1 U1424 ( .A(n487), .B(n506), .Y(n3195) );
  XOR2X1 U1425 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B(n502), .Y(n3247) );
  XOR2X1 U1426 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B(n477), .Y(n3255) );
  XOR2X1 U1427 ( .A(n491), .B(n511), .Y(n3215) );
  XOR2X1 U1428 ( .A(n458), .B(n486), .Y(n3205) );
  XOR2X1 U1429 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B(n468), .Y(n3257) );
  XOR2X1 U1430 ( .A(n450), .B(n476), .Y(n3209) );
  XOR2X1 U1431 ( .A(n435), .B(n434), .Y(n3265) );
  OR3XL U1432 ( .A(results_a1_a2[11]), .B(results_a1_a2[12]), 
        .C(results_a1_a2_inv_inverterxn15), .Y(results_a1_a2_inv_inverterxn13)
         );
  AND2X2 U1433 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer2_127827304_127827416)
         );
  AND2X2 U1434 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer2_127827752_127827920)
         );
  XOR2X1 U1435 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b8), .B(n3121), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831232_127845488_127847392)
         );
  XOR2X1 U1436 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b7), .B(n3137), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673456_127675360_127730576)
         );
  XOR2X1 U1437 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127827752_127827920)
         );
  XOR2X1 U1438 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .B(n3199), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128221424_128221536_128221704)
         );
  XOR2X1 U1439 ( .A(n467), .B(n3213), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127715424_128223048_128223272)
         );
  XNOR2X1 U1440 ( .A(n59), .B(results_a1_a2[4]), .Y(results_a1_a2_inv[4]) );
  NOR2X1 U1441 ( .A(results_a1_a2[3]), .B(results_a1_a2_inv_inverterxn8), 
        .Y(n59) );
  XNOR2X1 U1442 ( .A(n60), .B(results_a1_a2[6]), .Y(results_a1_a2_inv[6]) );
  NOR2X1 U1443 ( .A(results_a1_a2[5]), .B(results_a1_a2_inv_inverterxn6), 
        .Y(n60) );
  XNOR2X1 U1444 ( .A(n61), .B(results_a1_a2[8]), .Y(results_a1_a2_inv[8]) );
  NOR2X1 U1445 ( .A(results_a1_a2[7]), .B(results_a1_a2_inv_inverterxn4), 
        .Y(n61) );
  XOR2X1 U1446 ( .A(results_a1_a2_inv_inverterxn17), .B(results_a1_a2[10]), 
        .Y(results_a1_a2_inv[10]) );
  NAND2X1 U1447 ( .A(results_a1_a2_inv_inverterxn2), .B(n1302), 
        .Y(results_a1_a2_inv_inverterxn17) );
  XNOR2X1 U1448 ( .A(n62), .B(results_a1_a2[12]), .Y(results_a1_a2_inv[12]) );
  NOR2X1 U1449 ( .A(results_a1_a2_inv_inverterxn15), .B(results_a1_a2[11]), 
        .Y(n62) );
  XNOR2X1 U1450 ( .A(n63), .B(results_a1_a2[14]), .Y(results_a1_a2_inv[14]) );
  NOR2X1 U1451 ( .A(results_a1_a2[13]), .B(results_a1_a2_inv_inverterxn13), 
        .Y(n63) );
  XOR2X1 U1452 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b10), .B(n3135), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831456_127845712_127847616)
         );
  XOR2X1 U1453 ( .A(results_b0_b1_b2[16]), .B(results_a1_a2_inv[16]), 
        .Y(n4171) );
  XOR2X1 U1454 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127827304_127827416)
         );
  XOR2X1 U1455 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .B(n3195), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127827248_127827472_127827640)
         );
  XOR2X1 U1456 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .B(n3191), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127826576_127826800_127826968)
         );
  XOR2X1 U1457 ( 
        .A(output_p1_times_a1_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .B(n3197), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127827584_127827808_128221256)
         );
  XOR2X1 U1458 ( .A(n499), .B(n3209), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128222376_128222600_128222768)
         );
  OR3XL U1459 ( .A(results_a1_a2[3]), .B(results_a1_a2[4]), 
        .C(results_a1_a2_inv_inverterxn8), .Y(results_a1_a2_inv_inverterxn6)
         );
  XOR2X1 U1460 ( .A(n492), .B(n3201), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127635584_128221368_128221592)
         );
  XOR2X1 U1461 ( .A(n505), .B(n3205), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128221872_128222096_128222264)
         );
  XOR2X1 U1462 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .B(n3211), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128222936_128223104_128223216)
         );
  INVX1 U1463 ( .A(n4550), .Y(n480) );
  AOI22X1 U1464 ( .A0(n2353), .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[7]), 
        .B1(n4548), .Y(n4550) );
  XOR2X1 U1465 ( .A(n3809), .B(n2353), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[7]) );
  AND2X2 U1466 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n510), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer3_128246112_128246336)
         );
  BUFX3 U1467 ( .A(n4537), .Y(n229) );
  AOI22X1 U1468 ( .A0(\output_signal[2] ), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_2_), .B1(n165), 
        .Y(n4537) );
  XNOR2X1 U1469 ( .A(\output_signal[2] ), .B(n3782), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_2_) );
  NOR2XL U1470 ( .A(\output_signal[0] ), .B(\output_signal[1] ), .Y(n3782) );
  INVX1 U1471 ( .A(n4559), .Y(n408) );
  AOI22X1 U1472 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_15), 
        .A1(n113), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[15]), 
        .B1(n4548), .Y(n4559) );
  XNOR2X1 U1473 ( .A(n3817), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_15), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[15]) );
  INVX1 U1474 ( .A(n4549), .Y(n473) );
  AOI22X1 U1475 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_8), 
        .A1(n113), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[8]), 
        .B1(n4548), .Y(n4549) );
  XOR2X1 U1476 ( .A(n3808), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_8), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[8]) );
  OR2X2 U1477 ( .A(n2353), .B(n3809), .Y(n3808) );
  INVX1 U1478 ( .A(n4560), .Y(n417) );
  AOI22X1 U1479 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_14), 
        .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[14]), 
        .B1(n4548), .Y(n4560) );
  XOR2X1 U1480 ( .A(n3819), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_14), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[14]) );
  OR2X2 U1481 ( .A(output_p1_times_a1_mul_componentxunsigned_output_13), 
        .B(n3818), .Y(n3819) );
  BUFX3 U1482 ( .A(n4536), .Y(n228) );
  AOI22X1 U1483 ( .A0(\output_signal[3] ), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_3_), .B1(n165), 
        .Y(n4536) );
  XOR2X1 U1484 ( .A(n3781), .B(\output_signal[3] ), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_3_) );
  XOR2X1 U1485 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127672560_127674464), 
        .B(n3189), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127826464_127826632_127826744)
         );
  XOR2X1 U1486 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .B(n3187), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127672448_127826240_127826520)
         );
  XOR2X1 U1487 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .B(n3203), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128221760_128221928_128222040)
         );
  XOR2X1 U1488 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .B(n3207), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128222432_128222544_128222712)
         );
  XOR2X1 U1489 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n510), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128246112_128246336)
         );
  BUFX3 U1490 ( .A(n4535), .Y(n227) );
  AOI22X1 U1491 ( .A0(\output_signal[4] ), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_4_), .B1(n165), 
        .Y(n4535) );
  XOR2X1 U1492 ( .A(n3780), .B(\output_signal[4] ), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_4_) );
  OR2X2 U1493 ( .A(\output_signal[3] ), .B(n3781), .Y(n3780) );
  INVX1 U1494 ( .A(n4562), .Y(n432) );
  AOI22X1 U1495 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_12), 
        .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[12]), 
        .B1(n4548), .Y(n4562) );
  XOR2X1 U1496 ( .A(n3821), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_12), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[12]) );
  OR2X2 U1497 ( .A(n3820), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_11), .Y(n3821) );
  INVX1 U1498 ( .A(n4564), .Y(n453) );
  AOI22X1 U1499 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_10), 
        .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[10]), 
        .B1(n4548), .Y(n4564) );
  XOR2X1 U1500 ( .A(n3822), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_10), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[10]) );
  NAND2X1 U1501 ( .A(n3807), .B(n462), .Y(n3822) );
  BUFX3 U1502 ( .A(n4534), .Y(n226) );
  AOI22X1 U1503 ( .A0(\output_signal[5] ), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_5_), .B1(n165), 
        .Y(n4534) );
  XOR2X1 U1504 ( .A(n3779), .B(\output_signal[5] ), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_5_) );
  BUFX3 U1505 ( .A(n4533), .Y(n225) );
  AOI22X1 U1506 ( .A0(\output_signal[6] ), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_6_), .B1(n165), 
        .Y(n4533) );
  XOR2X1 U1507 ( .A(n3778), .B(\output_signal[6] ), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_6_) );
  OR2X2 U1508 ( .A(\output_signal[5] ), .B(n3779), .Y(n3778) );
  INVX1 U1509 ( .A(n3128), .Y(n436) );
  AOI22X1 U1510 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b10), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b11), .B0(n3127), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b9), .Y(n3128) );
  INVX1 U1511 ( .A(n3190), .Y(n502) );
  AOI22X1 U1512 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .A1(n508), .B0(n3189), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127672560_127674464), 
        .Y(n3190) );
  INVX1 U1513 ( .A(n3198), .Y(n477) );
  AOI22X1 U1514 ( .A0(n500), .A1(n479), .B0(n3197), 
        .B1(output_p1_times_a1_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .Y(n3198) );
  INVX1 U1515 ( .A(n3208), .Y(n451) );
  AOI22X1 U1516 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B0(n3207), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .Y(n3208) );
  INVX1 U1517 ( .A(n3212), .Y(n439) );
  AOI22X1 U1518 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .A1(output_p1_times_a1_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B0(n3211), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .Y(n3212) );
  INVX1 U1519 ( .A(n3266), .Y(n433) );
  AOI22X1 U1520 ( .A0(n434), .A1(n435), .B0(n3265), .B1(n456), .Y(n3266) );
  BUFX3 U1521 ( .A(n4532), .Y(n224) );
  AOI22X1 U1522 ( .A0(\output_signal[7] ), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_7_), .B1(n165), 
        .Y(n4532) );
  XOR2X1 U1523 ( .A(n3777), .B(\output_signal[7] ), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_7_) );
  INVX1 U1524 ( .A(n4563), .Y(n441) );
  AOI22X1 U1525 ( .A0(output_p1_times_a1_mul_componentxunsigned_output_11), 
        .A1(n113), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[11]), 
        .B1(n4548), .Y(n4563) );
  XOR2X1 U1526 ( .A(n3820), 
        .B(output_p1_times_a1_mul_componentxunsigned_output_11), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[11]) );
  INVX1 U1527 ( .A(n3196), .Y(n483) );
  AOI22X1 U1528 ( .A0(n506), .A1(n487), .B0(n3195), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .Y(n3196) );
  INVX1 U1529 ( .A(n3256), .Y(n470) );
  AOI22X1 U1530 ( .A0(n477), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B0(n3255), .B1(n471), .Y(n3256) );
  INVX1 U1531 ( .A(n3258), .Y(n459) );
  AOI22X1 U1532 ( .A0(n468), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B0(n3257), .B1(n461), .Y(n3258) );
  INVX1 U1533 ( .A(n3210), .Y(n447) );
  AOI22X1 U1534 ( .A0(n476), .A1(n450), .B0(n3209), .B1(n499), .Y(n3210) );
  BUFX3 U1535 ( .A(n4531), .Y(n223) );
  AOI22X1 U1536 ( .A0(output_previous_1[8]), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_8_), .B1(n165), 
        .Y(n4531) );
  XOR2X1 U1537 ( .A(n3776), .B(output_previous_1[8]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_8_) );
  OR2X2 U1538 ( .A(\output_signal[7] ), .B(n3777), .Y(n3776) );
  INVX1 U1539 ( .A(n3200), .Y(n471) );
  AOI22X1 U1540 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B0(n3199), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .Y(n3200) );
  INVX1 U1541 ( .A(n3248), .Y(n496) );
  AOI22X1 U1542 ( .A0(n502), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B0(n3247), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .Y(n3248) );
  BUFX3 U1543 ( .A(n4530), .Y(n222) );
  AOI22X1 U1544 ( .A0(output_previous_1[9]), .A1(n134), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_9_), .B1(n165), 
        .Y(n4530) );
  XNOR2X1 U1545 ( .A(n3775), .B(output_previous_1[9]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_9_) );
  INVX1 U1546 ( .A(results_a1_a2[9]), .Y(n1302) );
  AOI22X1 U1547 ( .A0(output_previous_1[12]), .A1(n133), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_12_), .B1(n165), 
        .Y(n4543) );
  XOR2X1 U1548 ( .A(n3789), .B(output_previous_1[12]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_12_) );
  OR2X2 U1549 ( .A(n3788), .B(output_previous_1[11]), .Y(n3789) );
  AOI22X1 U1550 ( .A0(output_previous_1[13]), .A1(n133), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_13_), .B1(n165), 
        .Y(n4542) );
  XOR2X1 U1551 ( .A(n3786), .B(output_previous_1[13]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_13_) );
  INVX1 U1552 ( .A(n3136), .Y(n428) );
  AOI22X1 U1553 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b11), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b12), .B0(n3135), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b10), .Y(n3136) );
  INVX1 U1554 ( .A(n3146), .Y(n446) );
  AOI22X1 U1555 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b9), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b10), .B0(n3145), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b8), .Y(n3146) );
  INVX1 U1556 ( .A(n3144), .Y(n426) );
  AOI22X1 U1557 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b12), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b13), .B0(n3143), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b11), .Y(n3144) );
  INVX1 U1558 ( .A(n4552), .Y(n495) );
  AOI22X1 U1559 ( .A0(output_p1_times_a1_mul_componentxUMxfirst_vector[5]), 
        .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[5]), 
        .B1(n4548), .Y(n4552) );
  XOR2X1 U1560 ( .A(n3811), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[5]), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[5]) );
  INVX1 U1561 ( .A(n3228), .Y(n442) );
  AOI22X1 U1562 ( 
        .A0(output_p1_times_a1_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .A1(n498), .B0(n3227), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .Y(n3228) );
  AOI22X1 U1563 ( .A0(n507), .A1(n484), .B0(n3239), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .Y(n3240) );
  INVX1 U1564 ( .A(n3138), .Y(n455) );
  AOI22X1 U1565 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b8), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b9), .B0(n3137), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b7), .Y(n3138) );
  INVX1 U1566 ( .A(n3234), .Y(n465) );
  AOI22X1 U1567 ( .A0(n490), .A1(n466), .B0(n3233), .B1(n514), .Y(n3234) );
  OR3XL U1568 ( .A(\output_signal[1] ), .B(\output_signal[2] ), 
        .C(\output_signal[0] ), .Y(n3781) );
  XOR2X1 U1569 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[2]) );
  XOR2X1 U1570 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b10), .B(n3163), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673792_127675696_127730912)
         );
  XOR2X1 U1571 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b10), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b9), .Y(n3145) );
  XOR2X1 U1572 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b11), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b10), .Y(n3153) );
  XOR2X1 U1573 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b12), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b11), .Y(n3163) );
  XOR2X1 U1574 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b14), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b13), .Y(n3151) );
  XOR2X1 U1575 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b15), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b14), .Y(n3161) );
  XOR2X1 U1576 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b8), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b7), .Y(n3155) );
  XOR2X1 U1577 ( .A(n474), .B(n3225), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128224392_128224616_128224784)
         );
  XOR2X1 U1578 ( .A(n514), .B(n3233), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128197016_128197240_128197352)
         );
  XOR2X1 U1579 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .Y(n3223) );
  XOR2X1 U1580 ( .A(n498), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .Y(n3227) );
  XOR2X1 U1581 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .Y(n3229) );
  XOR2X1 U1582 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B(n427), .Y(n3269) );
  XOR2X1 U1583 ( .A(n466), .B(n490), .Y(n3233) );
  XOR2X1 U1584 ( .A(n484), .B(n507), .Y(n3239) );
  XOR2X1 U1585 ( .A(n410), .B(n465), .Y(n3277) );
  XOR2X1 U1586 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b13), .B(n3161), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831792_127846048_127847952)
         );
  XOR2X1 U1587 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b9), .B(n3153), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673680_127675584_127730800)
         );
  XOR2X1 U1588 ( .A(n485), .B(n3219), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128223720_128223944_128224168)
         );
  XOR2X1 U1589 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .B(n3229), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128196792_128196960_128197184)
         );
  XOR2X1 U1590 ( .A(n411), .B(n3231), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_127627392_128196680_128196848)
         );
  XOR2X1 U1591 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b12), .B(n3151), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831680_127845936_127847840)
         );
  XOR2X1 U1592 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b8), .B(n3145), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673568_127675472_127730688)
         );
  XOR2X1 U1593 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .B(n3217), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128223888_128224112_128224056)
         );
  XOR2X1 U1594 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127715536_127848576), 
        .B(n3223), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128224728_128224896_128225064)
         );
  OR3XL U1595 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[3]), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[4]), .C(n3813), 
        .Y(n3811) );
  AND2X2 U1596 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer2_128223384_128223552)
         );
  AND2X2 U1597 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(output_p1_times_a1_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer2_127826128_127826296)
         );
  XOR2X1 U1598 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128263336_128263560_128263728), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer3_128263896_128264064_128264176), 
        .Y(n3304) );
  XOR2X1 U1599 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128198864_128199032_128199200), 
        .B(n3282), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128263896_128264064_128264176)
         );
  XOR2X1 U1600 ( .A(n399), .B(n3281), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128263336_128263560_128263728)
         );
  XOR2X1 U1601 ( 
        .A(output_p1_times_a1_mul_componentxUMxcarry_layer1_127627504_127629408), 
        .B(n3244), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128198864_128199032_128199200)
         );
  XOR2X1 U1602 ( .A(n400), 
        .B(output_p1_times_a1_mul_componentxUMxsecond_vector[17]), .Y(n2355)
         );
  XOR2X1 U1603 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer5_128315744_128315968_128316136), 
        .B(n3324), .Y(output_p1_times_a1_mul_componentxUMxsecond_vector[17])
         );
  INVX1 U1604 ( .A(n3323), .Y(n400) );
  XOR2X1 U1605 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128237752_128237976_128238144), 
        .B(n3319), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer5_128315744_128315968_128316136)
         );
  XOR2X1 U1606 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128223384_128223552)
         );
  INVX1 U1607 ( .A(n4553), .Y(n503) );
  AOI22X1 U1608 ( .A0(output_p1_times_a1_mul_componentxUMxfirst_vector[4]), 
        .A1(n113), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[4]), 
        .B1(n4548), .Y(n4553) );
  XOR2X1 U1609 ( .A(n3812), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[4]), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[4]) );
  OR2X2 U1610 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[3]), 
        .B(n3813), .Y(n3812) );
  INVX1 U1611 ( .A(n4551), .Y(n488) );
  AOI22XL U1612 ( .A0(output_p1_times_a1_mul_componentxUMxfirst_vector[6]), 
        .A1(n113), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[6]), 
        .B1(n4548), .Y(n4551) );
  XOR2X1 U1613 ( .A(n3810), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[6]), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[6]) );
  OR2X2 U1614 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[5]), 
        .B(n3811), .Y(n3810) );
  INVX1 U1615 ( .A(n3164), .Y(n403) );
  AOI22X1 U1616 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b11), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b12), .B0(n3163), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b10), .Y(n3164) );
  INVX1 U1617 ( .A(n3152), .Y(n443) );
  AOI22X1 U1618 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b13), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b14), .B0(n3151), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b12), .Y(n3152) );
  INVX1 U1619 ( .A(n3220), .Y(n427) );
  AOI22X1 U1620 ( .A0(n455), .A1(n428), .B0(n3219), .B1(n485), .Y(n3220) );
  INVX1 U1621 ( .A(n3270), .Y(n419) );
  AOI22X1 U1622 ( .A0(n427), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B0(n3269), .B1(n420), .Y(n3270) );
  AOI22X1 U1623 ( .A0(output_previous_1[14]), .A1(n133), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_14_), .B1(n165), 
        .Y(n4541) );
  XOR2X1 U1624 ( .A(n3787), .B(output_previous_1[14]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_14_) );
  OR2X2 U1625 ( .A(output_previous_1[13]), .B(n3786), .Y(n3787) );
  INVX1 U1626 ( .A(n3162), .Y(n444) );
  AOI22X1 U1627 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b14), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b15), .B0(n3161), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b13), .Y(n3162) );
  INVX1 U1628 ( .A(n3224), .Y(n475) );
  AOI22X1 U1629 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B0(n3223), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127715536_127848576), 
        .Y(n3224) );
  INVX1 U1630 ( .A(n3226), .Y(n424) );
  AOI22X1 U1631 ( .A0(n446), .A1(n426), .B0(n3225), .B1(n474), .Y(n3226) );
  INVX1 U1632 ( .A(n3154), .Y(n411) );
  AOI22X1 U1633 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b10), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b11), .B0(n3153), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b9), .Y(n3154) );
  INVX1 U1634 ( .A(n3222), .Y(n420) );
  AOI22X1 U1635 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .A1(n504), .B0(n3221), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .Y(n3222) );
  INVX1 U1636 ( .A(n3230), .Y(n413) );
  AOI22X1 U1637 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B0(n3229), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .Y(n3230) );
  AOI22X1 U1638 ( .A0(output_previous_1[15]), .A1(n133), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_15_), .B1(n165), 
        .Y(n4540) );
  XNOR2X1 U1639 ( .A(n3785), .B(output_previous_1[15]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_15_) );
  AOI22X1 U1640 ( .A0(output_previous_1[16]), .A1(n133), 
        .B0(output_p1_times_a1_mul_componentxinput_A_inverted_16_), .B1(n165), 
        .Y(n4539) );
  XNOR2X1 U1641 ( .A(n3784), .B(output_previous_1[16]), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_16_) );
  AOI22X1 U1642 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b9), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b10), .B0(n3175), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b8), .Y(n3176) );
  AOI22X1 U1643 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b12), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b13), .B0(n3173), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b11), .Y(n3174) );
  XOR2X1 U1644 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b8), .B(n3175), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732928_127722608_127724512)
         );
  XOR2X1 U1645 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b10), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b9), .Y(n3175) );
  XOR2X1 U1646 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b13), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b12), .Y(n3173) );
  XOR2X1 U1647 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b16), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b15), .Y(n3171) );
  XOR2X1 U1648 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b9), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b8), .Y(n3165) );
  XOR2X1 U1649 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b11), .B(n3173), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673904_127675808_127731024)
         );
  XOR2X1 U1650 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128198024_128197968)
         );
  XOR2X1 U1651 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b14), .B(n3171), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831904_127846160_127848064)
         );
  XOR2X1 U1652 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b7), .B(n3165), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732816_127722496_127724400)
         );
  OR3XL U1653 ( .A(n517), .B(n516), .C(n518), .Y(n4003) );
  XOR2X1 U1654 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .B(n3241), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128198472_128198640_128198808)
         );
  AND2X2 U1655 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer2_128198024_128197968)
         );
  INVX1 U1656 ( .A(n4554), .Y(n509) );
  AOI22XL U1657 ( .A0(output_p1_times_a1_mul_componentxUMxfirst_vector[3]), 
        .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[3]), 
        .B1(n4548), .Y(n4554) );
  XOR2X1 U1658 ( .A(n3813), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[3]), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[3]) );
  XOR2X1 U1659 ( 
        .A(output_p1_times_a1_mul_componentxUMxcarry_layer2_128198976_128199144), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128198304_128198528_128198696), 
        .Y(n3282) );
  AND2X2 U1660 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer2_128198976_128199144)
         );
  XOR2X1 U1661 ( .A(n445), .B(n3243), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128198304_128198528_128198696)
         );
  INVX1 U1662 ( .A(n3176), .Y(n445) );
  XOR2X1 U1663 ( .A(n3172), .B(n3174), .Y(n3243) );
  AOI22X1 U1664 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b15), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b16), .B0(n3171), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b14), .Y(n3172) );
  XOR2X1 U1665 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128198976_128199144)
         );
  INVX1 U1666 ( .A(n3166), .Y(n454) );
  AOI22X1 U1667 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b8), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b9), .B0(n3165), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b7), .Y(n3166) );
  INVX1 U1668 ( .A(n3242), .Y(n399) );
  AOI22X1 U1669 ( 
        .A0(output_p1_times_a1_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .A1(output_p1_times_a1_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B0(n3241), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .Y(n3242) );
  INVX1 U1670 ( .A(n3278), .Y(n404) );
  AOI22X1 U1671 ( .A0(n465), .A1(n410), .B0(n3277), .B1(n406), .Y(n3278) );
  XOR2X1 U1672 ( .A(n3783), .B(n165), 
        .Y(output_p1_times_a1_mul_componentxinput_A_inverted_17_) );
  NAND2BX1 U1673 ( .AN(output_previous_1[16]), .B(n3784), .Y(n3783) );
  XNOR2X1 U1674 ( .A(n516), .B(n4004), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[2]) );
  NOR2X1 U1675 ( .A(n518), .B(n517), .Y(n4004) );
  INVX1 U1676 ( .A(n3032), .Y(n1068) );
  AOI22X1 U1677 ( .A0(n1069), .A1(n1070), .B0(n3031), .B1(n1092), .Y(n3032) );
  INVX1 U1678 ( .A(n3500), .Y(n591) );
  AOI22X1 U1679 ( .A0(n592), .A1(n593), .B0(n3499), .B1(n615), .Y(n3500) );
  XOR2X1 U1680 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .B(n2747), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128223440_128223608_128223776)
         );
  XOR2X1 U1681 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .B(n2981), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128223440_128223608_128223776)
         );
  XOR2X1 U1682 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .B(n3449), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128223440_128223608_128223776)
         );
  XOR2X1 U1683 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .B(n2513), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128223440_128223608_128223776)
         );
  XOR2X1 U1684 ( .A(n968), .B(n988), .Y(n2747) );
  XOR2X1 U1685 ( .A(n1127), .B(n1147), .Y(n2981) );
  XOR2X1 U1686 ( .A(n650), .B(n670), .Y(n3449) );
  XOR2X1 U1687 ( .A(n809), .B(n829), .Y(n2513) );
  XOR2X1 U1688 ( .A(n911), .B(n910), .Y(n2797) );
  XOR2X1 U1689 ( .A(n1070), .B(n1069), .Y(n3031) );
  XOR2X1 U1690 ( .A(n593), .B(n592), .Y(n3499) );
  XOR2X1 U1691 ( .A(n752), .B(n751), .Y(n2563) );
  BUFX3 U1692 ( .A(n4451), .Y(n190) );
  AOI22X1 U1693 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_17), 
        .A1(n125), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[17]), 
        .B1(n4442), .Y(n4451) );
  XOR2X1 U1694 ( .A(n3719), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_17), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[17]) );
  XOR2X1 U1695 ( .A(n2312), .B(n2313), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_17) );
  BUFX3 U1696 ( .A(n4504), .Y(n211) );
  AOI22X1 U1697 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_17), 
        .A1(n129), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[17]), 
        .B1(n4495), .Y(n4504) );
  XOR2X1 U1698 ( .A(n3767), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_17), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[17]) );
  XOR2X1 U1699 ( .A(n2333), .B(n2334), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_17) );
  BUFX3 U1700 ( .A(n4610), .Y(n253) );
  AOI22X1 U1701 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_17), 
        .A1(n117), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[17]), 
        .B1(n4601), .Y(n4610) );
  XOR2X1 U1702 ( .A(n3863), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_17), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[17]) );
  XOR2X1 U1703 ( .A(n2375), .B(n2376), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_17) );
  BUFX3 U1704 ( .A(input_times_b0_mul_componentxn100), .Y(n281) );
  AOI22X1 U1705 ( .A0(input_times_b0_mul_componentxunsigned_output_17), 
        .A1(n121), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[17]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn100) );
  XOR2X1 U1706 ( .A(n3671), 
        .B(input_times_b0_mul_componentxunsigned_output_17), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[17]) );
  XOR2X1 U1707 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn474), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn475), 
        .Y(input_times_b0_mul_componentxunsigned_output_17) );
  INVX1 U1708 ( .A(n2748), .Y(n910) );
  AOI22X1 U1709 ( .A0(n988), .A1(n968), .B0(n2747), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .Y(n2748) );
  INVX1 U1710 ( .A(n2982), .Y(n1069) );
  AOI22X1 U1711 ( .A0(n1147), .A1(n1127), .B0(n2981), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .Y(n2982) );
  INVX1 U1712 ( .A(n3450), .Y(n592) );
  AOI22X1 U1713 ( .A0(n670), .A1(n650), .B0(n3449), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .Y(n3450) );
  INVX1 U1714 ( .A(n2514), .Y(n751) );
  AOI22X1 U1715 ( .A0(n829), .A1(n809), .B0(n2513), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127831456_127845712_127847616), 
        .Y(n2514) );
  INVX1 U1716 ( .A(n2798), .Y(n909) );
  AOI22X1 U1717 ( .A0(n910), .A1(n911), .B0(n2797), .B1(n933), .Y(n2798) );
  INVX1 U1718 ( .A(n2564), .Y(n750) );
  AOI22X1 U1719 ( .A0(n751), .A1(n752), .B0(n2563), .B1(n774), .Y(n2564) );
  XOR2X1 U1720 ( .A(n517), .B(n518), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[1]) );
  INVX1 U1721 ( .A(n4510), .Y(n1076) );
  AOI22X1 U1722 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_11), 
        .A1(n129), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[11]), 
        .B1(n4495), .Y(n4510) );
  XOR2X1 U1723 ( .A(n3772), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_11), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[11]) );
  INVX1 U1724 ( .A(n4616), .Y(n599) );
  AOI22X1 U1725 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_11), 
        .A1(n117), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[11]), 
        .B1(n4601), .Y(n4616) );
  XOR2X1 U1726 ( .A(n3868), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_11), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[11]) );
  INVX1 U1727 ( .A(n2722), .Y(n979) );
  AOI22X1 U1728 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .A1(n985), .B0(n2721), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127672560_127674464), 
        .Y(n2722) );
  INVX1 U1729 ( .A(n2956), .Y(n1138) );
  AOI22X1 U1730 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .A1(n1144), .B0(n2955), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127672560_127674464), 
        .Y(n2956) );
  INVX1 U1731 ( .A(n3424), .Y(n661) );
  AOI22X1 U1732 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .A1(n667), .B0(n3423), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127672560_127674464), 
        .Y(n3424) );
  INVX1 U1733 ( .A(n2488), .Y(n820) );
  AOI22X1 U1734 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .A1(n826), .B0(n2487), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127672560_127674464), 
        .Y(n2488) );
  INVX1 U1735 ( .A(n2974), .Y(n1087) );
  AOI22X1 U1736 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B0(n2973), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .Y(n2974) );
  INVX1 U1737 ( .A(n3442), .Y(n610) );
  AOI22X1 U1738 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B0(n3441), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .Y(n3442) );
  INVX1 U1739 ( .A(n2756), .Y(n952) );
  AOI22X1 U1740 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B0(n2755), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127715536_127848576), 
        .Y(n2756) );
  INVX1 U1741 ( .A(n2978), .Y(n1074) );
  AOI22X1 U1742 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .A1(input_p2_times_b2_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B0(n2977), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .Y(n2978) );
  INVX1 U1743 ( .A(n3446), .Y(n597) );
  AOI22X1 U1744 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .A1(output_p2_times_a2_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B0(n3445), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .Y(n3446) );
  INVX1 U1745 ( .A(n2522), .Y(n793) );
  AOI22X1 U1746 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B0(n2521), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127715536_127848576), 
        .Y(n2522) );
  AOI22X1 U1747 ( .A0(n984), .A1(n961), .B0(n2771), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .Y(n2772) );
  AOI22X1 U1748 ( .A0(n1143), .A1(n1120), .B0(n3005), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .Y(n3006) );
  AOI22X1 U1749 ( .A0(n666), .A1(n643), .B0(n3473), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .Y(n3474) );
  AOI22X1 U1750 ( .A0(n825), .A1(n802), .B0(n2537), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .Y(n2538) );
  INVX1 U1751 ( .A(n2738), .Y(n934) );
  AOI22X1 U1752 ( .A0(n963), .A1(n935), .B0(n2737), .B1(n982), .Y(n2738) );
  INVX1 U1753 ( .A(n2972), .Y(n1093) );
  AOI22X1 U1754 ( .A0(n1122), .A1(n1094), .B0(n2971), .B1(n1141), .Y(n2972) );
  INVX1 U1755 ( .A(n3440), .Y(n616) );
  AOI22X1 U1756 ( .A0(n645), .A1(n617), .B0(n3439), .B1(n664), .Y(n3440) );
  INVX1 U1757 ( .A(n2504), .Y(n775) );
  AOI22X1 U1758 ( .A0(n804), .A1(n776), .B0(n2503), .B1(n823), .Y(n2504) );
  INVX1 U1759 ( .A(n3022), .Y(n1106) );
  AOI22X1 U1760 ( .A0(n1113), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B0(n3021), .B1(n1107), .Y(n3022) );
  INVX1 U1761 ( .A(n3490), .Y(n629) );
  AOI22X1 U1762 ( .A0(n636), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B0(n3489), .B1(n630), .Y(n3490) );
  INVX1 U1763 ( .A(n2742), .Y(n924) );
  AOI22X1 U1764 ( .A0(n953), .A1(n927), .B0(n2741), .B1(n976), .Y(n2742) );
  INVX1 U1765 ( .A(n2508), .Y(n765) );
  AOI22X1 U1766 ( .A0(n794), .A1(n768), .B0(n2507), .B1(n817), .Y(n2508) );
  XOR2X1 U1767 ( .A(n990), .B(n2725), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127731808_127826912_127827136)
         );
  XOR2X1 U1768 ( .A(n1149), .B(n2959), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127731808_127826912_127827136)
         );
  XOR2X1 U1769 ( .A(n672), .B(n3427), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127731808_127826912_127827136)
         );
  XOR2X1 U1770 ( .A(n831), .B(n2491), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127731808_127826912_127827136)
         );
  XOR2X1 U1771 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .B(n2753), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128224280_128224448_128224560)
         );
  XOR2X1 U1772 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .B(n2987), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128224280_128224448_128224560)
         );
  XOR2X1 U1773 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .B(n3455), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128224280_128224448_128224560)
         );
  XOR2X1 U1774 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .B(n2519), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128224280_128224448_128224560)
         );
  XOR2X1 U1775 ( .A(n991), .B(n2765), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128197016_128197240_128197352)
         );
  XOR2X1 U1776 ( .A(n1150), .B(n2999), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128197016_128197240_128197352)
         );
  XOR2X1 U1777 ( .A(n673), .B(n3467), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128197016_128197240_128197352)
         );
  XOR2X1 U1778 ( .A(n832), .B(n2531), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128197016_128197240_128197352)
         );
  XOR2X1 U1779 ( .A(n978), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .Y(n2723) );
  XOR2X1 U1780 ( .A(n1137), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .Y(n2957) );
  XOR2X1 U1781 ( .A(n660), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .Y(n3425) );
  XOR2X1 U1782 ( .A(n819), 
        .B(input_times_b0_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .Y(n2489) );
  XOR2X1 U1783 ( .A(n985), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .Y(n2721) );
  XOR2X1 U1784 ( .A(n1144), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .Y(n2955) );
  XOR2X1 U1785 ( .A(n667), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .Y(n3423) );
  XOR2X1 U1786 ( .A(n826), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127830560_127844816_127846720), 
        .Y(n2487) );
  XOR2X1 U1787 ( .A(n970), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .Y(n2783) );
  XOR2X1 U1788 ( .A(n989), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .Y(n2735) );
  XOR2X1 U1789 ( .A(n1129), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .Y(n3017) );
  XOR2X1 U1790 ( .A(n1148), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .Y(n2969) );
  XOR2X1 U1791 ( .A(n652), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .Y(n3485) );
  XOR2X1 U1792 ( .A(n671), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .Y(n3437) );
  XOR2X1 U1793 ( .A(n811), 
        .B(input_times_b0_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .Y(n2549) );
  XOR2X1 U1794 ( .A(n830), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .Y(n2501) );
  XOR2X1 U1795 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .Y(n2731) );
  XOR2X1 U1796 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .Y(n2965) );
  XOR2X1 U1797 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .Y(n3433) );
  XOR2X1 U1798 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .Y(n2497) );
  XOR2X1 U1799 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .Y(n2739) );
  XOR2X1 U1800 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .Y(n2973) );
  XOR2X1 U1801 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .Y(n3441) );
  XOR2X1 U1802 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .Y(n2505) );
  XOR2X1 U1803 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .Y(n2749) );
  XOR2X1 U1804 ( .A(n981), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .Y(n2753) );
  XOR2X1 U1805 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .Y(n2755) );
  XOR2X1 U1806 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .Y(n2983) );
  XOR2X1 U1807 ( .A(n1140), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .Y(n2987) );
  XOR2X1 U1808 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .Y(n2989) );
  XOR2X1 U1809 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .Y(n3451) );
  XOR2X1 U1810 ( .A(n663), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .Y(n3455) );
  XOR2X1 U1811 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .Y(n3457) );
  XOR2X1 U1812 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .Y(n2515) );
  XOR2X1 U1813 ( .A(n822), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .Y(n2519) );
  XOR2X1 U1814 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .Y(n2521) );
  XOR2X1 U1815 ( 
        .A(input_p1_times_b1_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .Y(n2743) );
  XOR2X1 U1816 ( 
        .A(input_p2_times_b2_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .Y(n2977) );
  XOR2X1 U1817 ( 
        .A(output_p2_times_a2_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .Y(n3445) );
  XOR2X1 U1818 ( 
        .A(input_times_b0_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .Y(n2509) );
  XOR2X1 U1819 ( .A(n975), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .Y(n2759) );
  XOR2X1 U1820 ( .A(n1134), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .Y(n2993) );
  XOR2X1 U1821 ( .A(n657), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .Y(n3461) );
  XOR2X1 U1822 ( .A(n816), 
        .B(input_times_b0_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .Y(n2525) );
  XOR2X1 U1823 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .Y(n2761) );
  XOR2X1 U1824 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .Y(n2527) );
  XOR2X1 U1825 ( .A(n964), .B(n983), .Y(n2727) );
  XOR2X1 U1826 ( .A(n956), .B(n977), .Y(n2729) );
  XOR2X1 U1827 ( .A(n1123), .B(n1142), .Y(n2961) );
  XOR2X1 U1828 ( .A(n1115), .B(n1136), .Y(n2963) );
  XOR2X1 U1829 ( .A(n646), .B(n665), .Y(n3429) );
  XOR2X1 U1830 ( .A(n638), .B(n659), .Y(n3431) );
  XOR2X1 U1831 ( .A(n805), .B(n824), .Y(n2493) );
  XOR2X1 U1832 ( .A(n797), .B(n818), .Y(n2495) );
  XOR2X1 U1833 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B(n979), .Y(n2779) );
  XOR2X1 U1834 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B(n1138), .Y(n3013) );
  XOR2X1 U1835 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B(n661), .Y(n3481) );
  XOR2X1 U1836 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B(n820), .Y(n2545) );
  XOR2X1 U1837 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B(n945), .Y(n2789) );
  XOR2X1 U1838 ( .A(n935), .B(n963), .Y(n2737) );
  XOR2X1 U1839 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B(n954), .Y(n2787) );
  XOR2X1 U1840 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B(n1104), .Y(n3023) );
  XOR2X1 U1841 ( .A(n1094), .B(n1122), .Y(n2971) );
  XOR2X1 U1842 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B(n1113), .Y(n3021) );
  XOR2X1 U1843 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B(n627), .Y(n3491) );
  XOR2X1 U1844 ( .A(n617), .B(n645), .Y(n3439) );
  XOR2X1 U1845 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B(n636), .Y(n3489) );
  XOR2X1 U1846 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B(n786), .Y(n2555) );
  XOR2X1 U1847 ( .A(n776), .B(n804), .Y(n2503) );
  XOR2X1 U1848 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B(n795), .Y(n2553) );
  XOR2X1 U1849 ( .A(n927), .B(n953), .Y(n2741) );
  XOR2X1 U1850 ( .A(n1086), .B(n1112), .Y(n2975) );
  XOR2X1 U1851 ( .A(n609), .B(n635), .Y(n3443) );
  XOR2X1 U1852 ( .A(n768), .B(n794), .Y(n2507) );
  XOR2X1 U1853 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B(n903), .Y(n2801) );
  XOR2X1 U1854 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B(n1062), .Y(n3035) );
  XOR2X1 U1855 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B(n585), .Y(n3503) );
  XOR2X1 U1856 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B(n744), .Y(n2567) );
  XOR2X1 U1857 ( .A(n943), .B(n967), .Y(n2765) );
  XOR2X1 U1858 ( .A(n1102), .B(n1126), .Y(n2999) );
  XOR2X1 U1859 ( .A(n625), .B(n649), .Y(n3467) );
  XOR2X1 U1860 ( .A(n784), .B(n808), .Y(n2531) );
  XOR2X1 U1861 ( .A(n961), .B(n984), .Y(n2771) );
  XOR2X1 U1862 ( .A(n1120), .B(n1143), .Y(n3005) );
  XOR2X1 U1863 ( .A(n643), .B(n666), .Y(n3473) );
  XOR2X1 U1864 ( .A(n802), .B(n825), .Y(n2537) );
  AND2X2 U1865 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer2_127827304_127827416)
         );
  AND2X2 U1866 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer2_127827304_127827416)
         );
  AND2X2 U1867 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer2_127827304_127827416)
         );
  AND2X2 U1868 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer2_127827304_127827416)
         );
  AND2X2 U1869 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer2_127827752_127827920)
         );
  AND2X2 U1870 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer2_127827752_127827920)
         );
  AND2X2 U1871 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer2_127827752_127827920)
         );
  AND2X2 U1872 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer2_127827752_127827920)
         );
  XOR2X1 U1873 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127827752_127827920)
         );
  XOR2X1 U1874 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127827752_127827920) );
  XOR2X1 U1875 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .B(n2731), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128221424_128221536_128221704)
         );
  XOR2X1 U1876 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .B(n2965), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128221424_128221536_128221704)
         );
  XOR2X1 U1877 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .B(n3433), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128221424_128221536_128221704)
         );
  XOR2X1 U1878 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .B(n2497), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128221424_128221536_128221704)
         );
  XOR2X1 U1879 ( .A(n944), .B(n2745), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127715424_128223048_128223272)
         );
  XOR2X1 U1880 ( .A(n1103), .B(n2979), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127715424_128223048_128223272)
         );
  XOR2X1 U1881 ( .A(n626), .B(n3447), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127715424_128223048_128223272)
         );
  XOR2X1 U1882 ( .A(n785), .B(n2511), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127715424_128223048_128223272)
         );
  XOR2X1 U1883 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .B(n2761), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128196792_128196960_128197184)
         );
  XOR2X1 U1884 ( .A(n887), .B(n2763), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127627392_128196680_128196848)
         );
  XOR2X1 U1885 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .B(n2995), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128196792_128196960_128197184)
         );
  XOR2X1 U1886 ( .A(n1046), .B(n2997), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127627392_128196680_128196848)
         );
  XOR2X1 U1887 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .B(n3463), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128196792_128196960_128197184)
         );
  XOR2X1 U1888 ( .A(n569), .B(n3465), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127627392_128196680_128196848)
         );
  XOR2X1 U1889 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .B(n2527), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128196792_128196960_128197184)
         );
  XOR2X1 U1890 ( .A(n728), .B(n2529), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127627392_128196680_128196848)
         );
  XOR2X1 U1891 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127827304_127827416)
         );
  XOR2X1 U1892 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127827304_127827416)
         );
  XOR2X1 U1893 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127827304_127827416)
         );
  XOR2X1 U1894 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127672784_127674688_127729904), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127830784_127845040_127846944), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127827304_127827416) );
  XOR2X1 U1895 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .B(n2727), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127827248_127827472_127827640)
         );
  XOR2X1 U1896 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .B(n2961), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127827248_127827472_127827640)
         );
  XOR2X1 U1897 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .B(n3429), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127827248_127827472_127827640)
         );
  XOR2X1 U1898 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .B(n2493), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127827248_127827472_127827640)
         );
  XOR2X1 U1899 ( 
        .A(input_p1_times_b1_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .B(n2729), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127827584_127827808_128221256)
         );
  XOR2X1 U1900 ( 
        .A(input_p2_times_b2_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .B(n2963), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127827584_127827808_128221256)
         );
  XOR2X1 U1901 ( 
        .A(output_p2_times_a2_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .B(n3431), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127827584_127827808_128221256)
         );
  XOR2X1 U1902 ( 
        .A(input_times_b0_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .B(n2495), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127827584_127827808_128221256)
         );
  XOR2X1 U1903 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .B(n2749), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128223888_128224112_128224056)
         );
  XOR2X1 U1904 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .B(n2759), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128224952_128225120_128225232)
         );
  XOR2X1 U1905 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .B(n2983), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128223888_128224112_128224056)
         );
  XOR2X1 U1906 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .B(n2993), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128224952_128225120_128225232)
         );
  XOR2X1 U1907 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .B(n3451), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128223888_128224112_128224056)
         );
  XOR2X1 U1908 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .B(n3461), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128224952_128225120_128225232)
         );
  XOR2X1 U1909 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .B(n2515), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128223888_128224112_128224056)
         );
  XOR2X1 U1910 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .B(n2525), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128224952_128225120_128225232)
         );
  XOR2X1 U1911 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127715536_127848576), 
        .B(n2755), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128224728_128224896_128225064)
         );
  XOR2X1 U1912 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127715536_127848576), 
        .B(n2989), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128224728_128224896_128225064)
         );
  XOR2X1 U1913 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127715536_127848576), 
        .B(n3457), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128224728_128224896_128225064)
         );
  XOR2X1 U1914 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127715536_127848576), 
        .B(n2521), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128224728_128224896_128225064)
         );
  XOR2X1 U1915 ( .A(n982), .B(n2737), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128221872_128222096_128222264)
         );
  XOR2X1 U1916 ( .A(n969), .B(n2733), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127635584_128221368_128221592)
         );
  XOR2X1 U1917 ( .A(n1141), .B(n2971), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128221872_128222096_128222264)
         );
  XOR2X1 U1918 ( .A(n1128), .B(n2967), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127635584_128221368_128221592)
         );
  XOR2X1 U1919 ( .A(n664), .B(n3439), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128221872_128222096_128222264)
         );
  XOR2X1 U1920 ( .A(n651), .B(n3435), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127635584_128221368_128221592)
         );
  XOR2X1 U1921 ( .A(n823), .B(n2503), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128221872_128222096_128222264)
         );
  XOR2X1 U1922 ( .A(n810), .B(n2499), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127635584_128221368_128221592)
         );
  XOR2X1 U1923 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .B(n2743), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128222936_128223104_128223216)
         );
  XOR2X1 U1924 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .B(n2977), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128222936_128223104_128223216)
         );
  XOR2X1 U1925 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .B(n3445), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128222936_128223104_128223216)
         );
  XOR2X1 U1926 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .B(n2509), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128222936_128223104_128223216)
         );
  AND2X2 U1927 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer2_128223384_128223552)
         );
  AND2X2 U1928 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer2_128223384_128223552)
         );
  AND2X2 U1929 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer2_128223384_128223552)
         );
  AND2X2 U1930 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer2_128223384_128223552)
         );
  INVX1 U1931 ( .A(n4455), .Y(n899) );
  AOI22X1 U1932 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_13), 
        .A1(n125), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[13]), 
        .B1(n4442), .Y(n4455) );
  XOR2X1 U1933 ( .A(n3722), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_13), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[13]) );
  INVX1 U1934 ( .A(n4508), .Y(n1058) );
  AOI22X1 U1935 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_13), 
        .A1(n129), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[13]), 
        .B1(n4495), .Y(n4508) );
  XOR2X1 U1936 ( .A(n3770), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_13), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[13]) );
  INVX1 U1937 ( .A(n4614), .Y(n581) );
  AOI22X1 U1938 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_13), 
        .A1(n117), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[13]), 
        .B1(n4601), .Y(n4614) );
  XOR2X1 U1939 ( .A(n3866), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_13), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[13]) );
  INVX1 U1940 ( .A(input_times_b0_mul_componentxn104), .Y(n740) );
  AOI22X1 U1941 ( .A0(input_times_b0_mul_componentxunsigned_output_13), 
        .A1(n121), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[13]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn104) );
  XOR2X1 U1942 ( .A(n3674), 
        .B(input_times_b0_mul_componentxunsigned_output_13), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[13]) );
  INVX1 U1943 ( .A(n4453), .Y(n884) );
  AOI22X1 U1944 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_15), 
        .A1(n125), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[15]), 
        .B1(n4442), .Y(n4453) );
  XNOR2X1 U1945 ( .A(n3721), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_15), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[15]) );
  INVX1 U1946 ( .A(input_times_b0_mul_componentxn102), .Y(n725) );
  AOI22X1 U1947 ( .A0(input_times_b0_mul_componentxunsigned_output_15), 
        .A1(n121), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[15]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn102) );
  XNOR2X1 U1948 ( .A(n3673), 
        .B(input_times_b0_mul_componentxunsigned_output_15), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[15]) );
  INVX1 U1949 ( .A(n4454), .Y(n893) );
  AOI22X1 U1950 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_14), 
        .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[14]), 
        .B1(n4442), .Y(n4454) );
  XOR2X1 U1951 ( .A(n3723), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_14), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[14]) );
  OR2X2 U1952 ( .A(input_p1_times_b1_mul_componentxunsigned_output_13), 
        .B(n3722), .Y(n3723) );
  INVX1 U1953 ( .A(n4507), .Y(n1052) );
  AOI22X1 U1954 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_14), 
        .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[14]), 
        .B1(n4495), .Y(n4507) );
  XOR2X1 U1955 ( .A(n3771), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_14), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[14]) );
  OR2X2 U1956 ( .A(input_p2_times_b2_mul_componentxunsigned_output_13), 
        .B(n3770), .Y(n3771) );
  INVX1 U1957 ( .A(n4613), .Y(n575) );
  AOI22X1 U1958 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_14), 
        .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[14]), 
        .B1(n4601), .Y(n4613) );
  XOR2X1 U1959 ( .A(n3867), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_14), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[14]) );
  OR2X2 U1960 ( .A(output_p2_times_a2_mul_componentxunsigned_output_13), 
        .B(n3866), .Y(n3867) );
  INVX1 U1961 ( .A(input_times_b0_mul_componentxn103), .Y(n734) );
  AOI22X1 U1962 ( .A0(input_times_b0_mul_componentxunsigned_output_14), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[14]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn103) );
  XOR2X1 U1963 ( .A(n3675), 
        .B(input_times_b0_mul_componentxunsigned_output_14), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[14]) );
  OR2X2 U1964 ( .A(input_times_b0_mul_componentxunsigned_output_13), .B(n3674), 
        .Y(n3675) );
  XOR2X1 U1965 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128263336_128263560_128263728), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer3_128263896_128264064_128264176), 
        .Y(n2836) );
  XOR2X1 U1966 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128198864_128199032_128199200), 
        .B(n2814), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128263896_128264064_128264176)
         );
  XOR2X1 U1967 ( .A(n874), .B(n2813), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128263336_128263560_128263728)
         );
  XOR2X1 U1968 ( 
        .A(input_p1_times_b1_mul_componentxUMxcarry_layer1_127627504_127629408), 
        .B(n2776), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128198864_128199032_128199200)
         );
  XOR2X1 U1969 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128263336_128263560_128263728), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer3_128263896_128264064_128264176), 
        .Y(n3070) );
  XOR2X1 U1970 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128198864_128199032_128199200), 
        .B(n3048), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128263896_128264064_128264176)
         );
  XOR2X1 U1971 ( .A(n1033), .B(n3047), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128263336_128263560_128263728)
         );
  XOR2X1 U1972 ( 
        .A(input_p2_times_b2_mul_componentxUMxcarry_layer1_127627504_127629408), 
        .B(n3010), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128198864_128199032_128199200)
         );
  XOR2X1 U1973 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128263336_128263560_128263728), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer3_128263896_128264064_128264176), 
        .Y(n3538) );
  XOR2X1 U1974 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128198864_128199032_128199200), 
        .B(n3516), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128263896_128264064_128264176)
         );
  XOR2X1 U1975 ( .A(n556), .B(n3515), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128263336_128263560_128263728)
         );
  XOR2X1 U1976 ( 
        .A(output_p2_times_a2_mul_componentxUMxcarry_layer1_127627504_127629408), 
        .B(n3478), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128198864_128199032_128199200)
         );
  XOR2X1 U1977 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128263336_128263560_128263728), 
        .B(input_times_b0_mul_componentxUMxsum_layer3_128263896_128264064_128264176), 
        .Y(n2602) );
  XOR2X1 U1978 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128198864_128199032_128199200), 
        .B(n2580), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128263896_128264064_128264176)
         );
  XOR2X1 U1979 ( .A(n715), .B(n2579), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128263336_128263560_128263728)
         );
  XOR2X1 U1980 ( 
        .A(input_times_b0_mul_componentxUMxcarry_layer1_127627504_127629408), 
        .B(n2542), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128198864_128199032_128199200)
         );
  XOR2X1 U1981 ( .A(n2770), .B(n2772), .Y(n2813) );
  AOI22X1 U1982 ( .A0(n879), .A1(n920), .B0(n2769), .B1(n931), .Y(n2770) );
  XOR2X1 U1983 ( .A(n3004), .B(n3006), .Y(n3047) );
  AOI22X1 U1984 ( .A0(n1038), .A1(n1079), .B0(n3003), .B1(n1090), .Y(n3004) );
  XOR2X1 U1985 ( .A(n3472), .B(n3474), .Y(n3515) );
  AOI22X1 U1986 ( .A0(n561), .A1(n602), .B0(n3471), .B1(n613), .Y(n3472) );
  XOR2X1 U1987 ( .A(n2536), .B(n2538), .Y(n2579) );
  AOI22X1 U1988 ( .A0(n720), .A1(n761), .B0(n2535), .B1(n772), .Y(n2536) );
  XOR2X1 U1989 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer4_128238312_128238424_128238592), 
        .B(n881), .Y(n2856) );
  XOR2X1 U1990 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer3_128264344_128264512), 
        .B(n2836), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer4_128238312_128238424_128238592)
         );
  INVX1 U1991 ( .A(n2850), .Y(n881) );
  XOR2X1 U1992 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_128199816_128200040_128199984), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128199368_128199480_128199648), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128264344_128264512)
         );
  XOR2X1 U1993 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer4_128238312_128238424_128238592), 
        .B(n1040), .Y(n3090) );
  XOR2X1 U1994 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer3_128264344_128264512), 
        .B(n3070), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer4_128238312_128238424_128238592)
         );
  INVX1 U1995 ( .A(n3084), .Y(n1040) );
  XOR2X1 U1996 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_128199816_128200040_128199984), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128199368_128199480_128199648), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128264344_128264512)
         );
  XOR2X1 U1997 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer4_128238312_128238424_128238592), 
        .B(n563), .Y(n3558) );
  XOR2X1 U1998 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer3_128264344_128264512), 
        .B(n3538), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer4_128238312_128238424_128238592)
         );
  INVX1 U1999 ( .A(n3552), .Y(n563) );
  XOR2X1 U2000 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_128199816_128200040_128199984), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128199368_128199480_128199648), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128264344_128264512)
         );
  XOR2X1 U2001 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer4_128238312_128238424_128238592), 
        .B(n722), .Y(n2622) );
  XOR2X1 U2002 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer3_128264344_128264512), 
        .B(n2602), 
        .Y(input_times_b0_mul_componentxUMxsum_layer4_128238312_128238424_128238592)
         );
  INVX1 U2003 ( .A(n2616), .Y(n722) );
  XOR2X1 U2004 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_128199816_128200040_128199984), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128199368_128199480_128199648), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128264344_128264512) );
  XOR2X1 U2005 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128223384_128223552)
         );
  XOR2X1 U2006 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128223384_128223552)
         );
  XOR2X1 U2007 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128223384_128223552)
         );
  XOR2X1 U2008 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127635808_127637712_127713408), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127732368_127722048_127723952), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128223384_128223552) );
  XOR2X1 U2009 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .B(n2739), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128222432_128222544_128222712)
         );
  XOR2X1 U2010 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .B(n2735), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128221760_128221928_128222040)
         );
  XOR2X1 U2011 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .B(n2973), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128222432_128222544_128222712)
         );
  XOR2X1 U2012 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .B(n2969), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128221760_128221928_128222040)
         );
  XOR2X1 U2013 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .B(n3441), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128222432_128222544_128222712)
         );
  XOR2X1 U2014 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .B(n3437), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128221760_128221928_128222040)
         );
  XOR2X1 U2015 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .B(n2505), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128222432_128222544_128222712)
         );
  XOR2X1 U2016 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .B(n2501), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128221760_128221928_128222040)
         );
  INVX1 U2017 ( .A(n4456), .Y(n908) );
  AOI22X1 U2018 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_12), 
        .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[12]), 
        .B1(n4442), .Y(n4456) );
  XOR2X1 U2019 ( .A(n3725), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_12), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[12]) );
  OR2X2 U2020 ( .A(n3724), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_11), .Y(n3725) );
  INVX1 U2021 ( .A(n4509), .Y(n1067) );
  AOI22X1 U2022 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_12), 
        .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[12]), 
        .B1(n4495), .Y(n4509) );
  XOR2X1 U2023 ( .A(n3773), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_12), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[12]) );
  OR2X2 U2024 ( .A(n3772), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_11), .Y(n3773) );
  INVX1 U2025 ( .A(n4615), .Y(n590) );
  AOI22X1 U2026 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_12), 
        .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[12]), 
        .B1(n4601), .Y(n4615) );
  XOR2X1 U2027 ( .A(n3869), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_12), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[12]) );
  OR2X2 U2028 ( .A(n3868), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_11), .Y(n3869) );
  INVX1 U2029 ( .A(input_times_b0_mul_componentxn105), .Y(n749) );
  AOI22X1 U2030 ( .A0(input_times_b0_mul_componentxunsigned_output_12), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[12]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn105) );
  XOR2X1 U2031 ( .A(n3677), 
        .B(input_times_b0_mul_componentxunsigned_output_12), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[12]) );
  OR2X2 U2032 ( .A(n3676), .B(input_times_b0_mul_componentxunsigned_output_11), 
        .Y(n3677) );
  INVX1 U2033 ( .A(n4458), .Y(n930) );
  AOI22X1 U2034 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_10), 
        .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[10]), 
        .B1(n4442), .Y(n4458) );
  XOR2X1 U2035 ( .A(n3726), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_10), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[10]) );
  NAND2X1 U2036 ( .A(n3711), .B(n939), .Y(n3726) );
  INVX1 U2037 ( .A(n4511), .Y(n1089) );
  AOI22X1 U2038 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_10), 
        .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[10]), 
        .B1(n4495), .Y(n4511) );
  XOR2X1 U2039 ( .A(n3774), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_10), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[10]) );
  NAND2X1 U2040 ( .A(n3759), .B(n1098), .Y(n3774) );
  INVX1 U2041 ( .A(n4617), .Y(n612) );
  AOI22X1 U2042 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_10), 
        .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[10]), 
        .B1(n4601), .Y(n4617) );
  XOR2X1 U2043 ( .A(n3870), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_10), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[10]) );
  NAND2X1 U2044 ( .A(n3855), .B(n621), .Y(n3870) );
  INVX1 U2045 ( .A(input_times_b0_mul_componentxn107), .Y(n771) );
  AOI22X1 U2046 ( .A0(input_times_b0_mul_componentxunsigned_output_10), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[10]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn107) );
  XOR2X1 U2047 ( .A(n3678), 
        .B(input_times_b0_mul_componentxunsigned_output_10), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[10]) );
  NAND2X1 U2048 ( .A(n3663), .B(n780), .Y(n3678) );
  INVX1 U2049 ( .A(n4452), .Y(n876) );
  AOI22X1 U2050 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_16), 
        .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[16]), 
        .B1(n4442), .Y(n4452) );
  XNOR2X1 U2051 ( .A(n3720), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_16), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[16]) );
  INVX1 U2052 ( .A(input_times_b0_mul_componentxn101), .Y(n717) );
  AOI22X1 U2053 ( .A0(input_times_b0_mul_componentxunsigned_output_16), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[16]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn101) );
  XNOR2X1 U2054 ( .A(n3672), 
        .B(input_times_b0_mul_componentxunsigned_output_16), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[16]) );
  INVX1 U2055 ( .A(n2730), .Y(n954) );
  AOI22X1 U2056 ( .A0(n977), .A1(n956), .B0(n2729), 
        .B1(input_p1_times_b1_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .Y(n2730) );
  INVX1 U2057 ( .A(n2964), .Y(n1113) );
  AOI22X1 U2058 ( .A0(n1136), .A1(n1115), .B0(n2963), 
        .B1(input_p2_times_b2_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .Y(n2964) );
  INVX1 U2059 ( .A(n3432), .Y(n636) );
  AOI22X1 U2060 ( .A0(n659), .A1(n638), .B0(n3431), 
        .B1(output_p2_times_a2_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .Y(n3432) );
  INVX1 U2061 ( .A(n2496), .Y(n795) );
  AOI22X1 U2062 ( .A0(n818), .A1(n797), .B0(n2495), 
        .B1(input_times_b0_mul_componentxUMxcarry_layer1_127731920_127721600), 
        .Y(n2496) );
  INVX1 U2063 ( .A(n2784), .Y(n959) );
  AOI22X1 U2064 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .A1(n970), .B0(n2783), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .Y(n2784) );
  INVX1 U2065 ( .A(n3018), .Y(n1118) );
  AOI22X1 U2066 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .A1(n1129), .B0(n3017), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .Y(n3018) );
  INVX1 U2067 ( .A(n3486), .Y(n641) );
  AOI22X1 U2068 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .A1(n652), .B0(n3485), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .Y(n3486) );
  INVX1 U2069 ( .A(n2550), .Y(n800) );
  AOI22X1 U2070 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer2_127827304_127827416), 
        .A1(n811), .B0(n2549), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_127827248_127827472_127827640), 
        .Y(n2550) );
  INVX1 U2071 ( .A(n2740), .Y(n928) );
  AOI22X1 U2072 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B0(n2739), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .Y(n2740) );
  INVX1 U2073 ( .A(n2506), .Y(n769) );
  AOI22X1 U2074 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127673232_127675136_127730352), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127831232_127845488_127847392), 
        .B0(n2505), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127732256_127721936_127723840), 
        .Y(n2506) );
  INVX1 U2075 ( .A(n2744), .Y(n915) );
  AOI22X1 U2076 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .A1(input_p1_times_b1_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B0(n2743), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .Y(n2744) );
  INVX1 U2077 ( .A(n2510), .Y(n756) );
  AOI22X1 U2078 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127831344_127845600_127847504), 
        .A1(input_times_b0_mul_componentxUMxcarry_layer1_127635696_127637600), 
        .B0(n2509), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127673344_127675248_127730464), 
        .Y(n2510) );
  INVX1 U2079 ( .A(n2802), .Y(n895) );
  AOI22X1 U2080 ( .A0(n903), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B0(n2801), .B1(n896), .Y(n2802) );
  INVX1 U2081 ( .A(n2760), .Y(n918) );
  AOI22X1 U2082 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .A1(n975), .B0(n2759), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .Y(n2760) );
  INVX1 U2083 ( .A(n3036), .Y(n1054) );
  AOI22X1 U2084 ( .A0(n1062), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B0(n3035), .B1(n1055), .Y(n3036) );
  INVX1 U2085 ( .A(n2994), .Y(n1077) );
  AOI22X1 U2086 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .A1(n1134), .B0(n2993), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .Y(n2994) );
  INVX1 U2087 ( .A(n3504), .Y(n577) );
  AOI22X1 U2088 ( .A0(n585), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B0(n3503), .B1(n578), .Y(n3504) );
  INVX1 U2089 ( .A(n3462), .Y(n600) );
  AOI22X1 U2090 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .A1(n657), .B0(n3461), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .Y(n3462) );
  INVX1 U2091 ( .A(n2568), .Y(n736) );
  AOI22X1 U2092 ( .A0(n744), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127715648_127848688_127850592), 
        .B0(n2567), .B1(n737), .Y(n2568) );
  INVX1 U2093 ( .A(n2526), .Y(n759) );
  AOI22X1 U2094 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer1_127715536_127848576), 
        .A1(n816), .B0(n2525), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127831680_127845936_127847840), 
        .Y(n2526) );
  INVX1 U2095 ( .A(n4506), .Y(n1043) );
  AOI22X1 U2096 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_15), 
        .A1(n129), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[15]), 
        .B1(n4495), .Y(n4506) );
  XNOR2X1 U2097 ( .A(n3769), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_15), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[15]) );
  INVX1 U2098 ( .A(n4612), .Y(n566) );
  AOI22X1 U2099 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_15), 
        .A1(n117), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[15]), 
        .B1(n4601), .Y(n4612) );
  XNOR2X1 U2100 ( .A(n3865), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_15), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[15]) );
  INVX1 U2101 ( .A(n4505), .Y(n1035) );
  AOI22X1 U2102 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_16), 
        .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[16]), 
        .B1(n4495), .Y(n4505) );
  XNOR2X1 U2103 ( .A(n3768), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_16), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[16]) );
  INVX1 U2104 ( .A(n4611), .Y(n558) );
  AOI22X1 U2105 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_16), 
        .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[16]), 
        .B1(n4601), .Y(n4611) );
  XNOR2X1 U2106 ( .A(n3864), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_16), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[16]) );
  INVX1 U2107 ( .A(n4457), .Y(n917) );
  AOI22X1 U2108 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_11), 
        .A1(n125), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[11]), 
        .B1(n4442), .Y(n4457) );
  XOR2X1 U2109 ( .A(n3724), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_11), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[11]) );
  INVX1 U2110 ( .A(input_times_b0_mul_componentxn106), .Y(n758) );
  AOI22X1 U2111 ( .A0(input_times_b0_mul_componentxunsigned_output_11), 
        .A1(n121), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[11]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn106) );
  XOR2X1 U2112 ( .A(n3676), 
        .B(input_times_b0_mul_componentxunsigned_output_11), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[11]) );
  BUFX3 U2113 ( .A(n254), .Y(n144) );
  BUFX3 U2114 ( .A(n282), .Y(n132) );
  INVX1 U2115 ( .A(n2724), .Y(n974) );
  AOI22X1 U2116 ( 
        .A0(input_p1_times_b1_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .A1(n978), .B0(n2723), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .Y(n2724) );
  INVX1 U2117 ( .A(n2958), .Y(n1133) );
  AOI22X1 U2118 ( 
        .A0(input_p2_times_b2_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .A1(n1137), .B0(n2957), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .Y(n2958) );
  INVX1 U2119 ( .A(n3426), .Y(n656) );
  AOI22X1 U2120 ( 
        .A0(output_p2_times_a2_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .A1(n660), .B0(n3425), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .Y(n3426) );
  INVX1 U2121 ( .A(n2490), .Y(n815) );
  AOI22X1 U2122 ( 
        .A0(input_times_b0_mul_componentxUMxcarry_layer1_127672560_127674464), 
        .A1(n819), .B0(n2489), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .Y(n2490) );
  INVX1 U2123 ( .A(n2728), .Y(n960) );
  AOI22X1 U2124 ( .A0(n983), .A1(n964), .B0(n2727), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .Y(n2728) );
  INVX1 U2125 ( .A(n2962), .Y(n1119) );
  AOI22X1 U2126 ( .A0(n1142), .A1(n1123), .B0(n2961), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .Y(n2962) );
  INVX1 U2127 ( .A(n3430), .Y(n642) );
  AOI22X1 U2128 ( .A0(n665), .A1(n646), .B0(n3429), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .Y(n3430) );
  INVX1 U2129 ( .A(n2494), .Y(n801) );
  AOI22X1 U2130 ( .A0(n824), .A1(n805), .B0(n2493), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127830896_127845152_127847056), 
        .Y(n2494) );
  INVX1 U2131 ( .A(n2790), .Y(n936) );
  AOI22X1 U2132 ( .A0(n945), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B0(n2789), .B1(n938), .Y(n2790) );
  INVX1 U2133 ( .A(n2788), .Y(n947) );
  AOI22X1 U2134 ( .A0(n954), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B0(n2787), .B1(n948), .Y(n2788) );
  INVX1 U2135 ( .A(n3024), .Y(n1095) );
  AOI22X1 U2136 ( .A0(n1104), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B0(n3023), .B1(n1097), .Y(n3024) );
  INVX1 U2137 ( .A(n3492), .Y(n618) );
  AOI22X1 U2138 ( .A0(n627), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B0(n3491), .B1(n620), .Y(n3492) );
  INVX1 U2139 ( .A(n2556), .Y(n777) );
  AOI22X1 U2140 ( .A0(n786), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127635696_127637600), 
        .B0(n2555), .B1(n779), .Y(n2556) );
  INVX1 U2141 ( .A(n2554), .Y(n788) );
  AOI22X1 U2142 ( .A0(n795), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127732144_127721824_127723728), 
        .B0(n2553), .B1(n789), .Y(n2554) );
  INVX1 U2143 ( .A(n2976), .Y(n1083) );
  AOI22X1 U2144 ( .A0(n1112), .A1(n1086), .B0(n2975), .B1(n1135), .Y(n2976) );
  INVX1 U2145 ( .A(n2990), .Y(n1111) );
  AOI22X1 U2146 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B0(n2989), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127715536_127848576), 
        .Y(n2990) );
  INVX1 U2147 ( .A(n3444), .Y(n606) );
  AOI22X1 U2148 ( .A0(n635), .A1(n609), .B0(n3443), .B1(n658), .Y(n3444) );
  INVX1 U2149 ( .A(n3458), .Y(n634) );
  AOI22X1 U2150 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127636032_127637936_127713632), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127732592_127722272_127724176), 
        .B0(n3457), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127715536_127848576), 
        .Y(n3458) );
  INVX1 U2151 ( .A(n2736), .Y(n938) );
  AOI22X1 U2152 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .A1(n989), .B0(n2735), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .Y(n2736) );
  INVX1 U2153 ( .A(n2732), .Y(n948) );
  AOI22X1 U2154 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B0(n2731), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .Y(n2732) );
  INVX1 U2155 ( .A(n2970), .Y(n1097) );
  AOI22X1 U2156 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .A1(n1148), .B0(n2969), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .Y(n2970) );
  INVX1 U2157 ( .A(n2966), .Y(n1107) );
  AOI22X1 U2158 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B0(n2965), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .Y(n2966) );
  INVX1 U2159 ( .A(n3438), .Y(n620) );
  AOI22X1 U2160 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .A1(n671), .B0(n3437), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .Y(n3438) );
  INVX1 U2161 ( .A(n3434), .Y(n630) );
  AOI22X1 U2162 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B0(n3433), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .Y(n3434) );
  INVX1 U2163 ( .A(n2502), .Y(n779) );
  AOI22X1 U2164 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127831120_127845376_127847280), 
        .A1(n830), .B0(n2501), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127673120_127675024_127730240), 
        .Y(n2502) );
  INVX1 U2165 ( .A(n2498), .Y(n789) );
  AOI22X1 U2166 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127673008_127674912_127730128), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127831008_127845264_127847168), 
        .B0(n2497), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127732032_127721712_127723616), 
        .Y(n2498) );
  INVX1 U2167 ( .A(n2750), .Y(n933) );
  AOI22X1 U2168 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B0(n2749), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .Y(n2750) );
  INVX1 U2169 ( .A(n2754), .Y(n896) );
  AOI22X1 U2170 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .A1(n981), .B0(n2753), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .Y(n2754) );
  INVX1 U2171 ( .A(n2984), .Y(n1092) );
  AOI22X1 U2172 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B0(n2983), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .Y(n2984) );
  INVX1 U2173 ( .A(n2988), .Y(n1055) );
  AOI22X1 U2174 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .A1(n1140), .B0(n2987), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .Y(n2988) );
  INVX1 U2175 ( .A(n3452), .Y(n615) );
  AOI22X1 U2176 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B0(n3451), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .Y(n3452) );
  INVX1 U2177 ( .A(n3456), .Y(n578) );
  AOI22X1 U2178 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .A1(n663), .B0(n3455), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .Y(n3456) );
  INVX1 U2179 ( .A(n2516), .Y(n774) );
  AOI22X1 U2180 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127732480_127722160_127724064), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127673456_127675360_127730576), 
        .B0(n2515), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127635920_127637824_127713520), 
        .Y(n2516) );
  INVX1 U2181 ( .A(n2520), .Y(n737) );
  AOI22X1 U2182 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127831568_127845824_127847728), 
        .A1(n822), .B0(n2519), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127673568_127675472_127730688), 
        .Y(n2520) );
  INVX1 U2183 ( .A(n2780), .Y(n973) );
  AOI22X1 U2184 ( .A0(n979), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B0(n2779), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .Y(n2780) );
  INVX1 U2185 ( .A(n3014), .Y(n1132) );
  AOI22X1 U2186 ( .A0(n1138), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B0(n3013), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .Y(n3014) );
  INVX1 U2187 ( .A(n3482), .Y(n655) );
  AOI22X1 U2188 ( .A0(n661), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B0(n3481), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .Y(n3482) );
  INVX1 U2189 ( .A(n2546), .Y(n814) );
  AOI22X1 U2190 ( .A0(n820), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127672672_127674576_127729792), 
        .B0(n2545), 
        .B1(input_times_b0_mul_componentxUMxsum_layer2_127826576_127826800_127826968), 
        .Y(n2546) );
  BUFX3 U2191 ( .A(n254), .Y(n143) );
  BUFX3 U2192 ( .A(n282), .Y(n131) );
  BUFX3 U2193 ( .A(n255), .Y(n141) );
  BUFX3 U2194 ( .A(n256), .Y(n139) );
  BUFX3 U2195 ( .A(n255), .Y(n142) );
  BUFX3 U2196 ( .A(n256), .Y(n140) );
  AOI22X1 U2197 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_9), 
        .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[9]), 
        .B1(n4442), .Y(n4441) );
  XNOR2X1 U2198 ( .A(n3711), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_9), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[9]) );
  AOI22X1 U2199 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_9), 
        .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[9]), 
        .B1(n4495), .Y(n4494) );
  XNOR2X1 U2200 ( .A(n3759), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_9), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[9]) );
  AOI22X1 U2201 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_9), 
        .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[9]), 
        .B1(n4601), .Y(n4600) );
  XNOR2X1 U2202 ( .A(n3855), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_9), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[9]) );
  AOI22X1 U2203 ( .A0(input_times_b0_mul_componentxunsigned_output_9), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[9]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn90) );
  XNOR2X1 U2204 ( .A(n3663), 
        .B(input_times_b0_mul_componentxunsigned_output_9), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[9]) );
  INVX1 U2205 ( .A(n4497), .Y(n1116) );
  AOI22X1 U2206 ( .A0(n2332), .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[7]), 
        .B1(n4495), .Y(n4497) );
  XOR2X1 U2207 ( .A(n3761), .B(n2332), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[7]) );
  INVX1 U2208 ( .A(n4603), .Y(n639) );
  AOI22X1 U2209 ( .A0(n2374), .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[7]), 
        .B1(n4601), .Y(n4603) );
  XOR2X1 U2210 ( .A(n3857), .B(n2374), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[7]) );
  INVX1 U2211 ( .A(n3008), .Y(n1033) );
  AOI22X1 U2212 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B0(n3007), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .Y(n3008) );
  INVX1 U2213 ( .A(n3476), .Y(n556) );
  AOI22X1 U2214 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B0(n3475), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .Y(n3476) );
  INVX1 U2215 ( .A(n2758), .Y(n900) );
  AOI22X1 U2216 ( .A0(n923), .A1(n902), .B0(n2757), .B1(n951), .Y(n2758) );
  INVX1 U2217 ( .A(n2992), .Y(n1059) );
  AOI22X1 U2218 ( .A0(n1082), .A1(n1061), .B0(n2991), .B1(n1110), .Y(n2992) );
  INVX1 U2219 ( .A(n3460), .Y(n582) );
  AOI22X1 U2220 ( .A0(n605), .A1(n584), .B0(n3459), .B1(n633), .Y(n3460) );
  INVX1 U2221 ( .A(n2524), .Y(n741) );
  AOI22X1 U2222 ( .A0(n764), .A1(n743), .B0(n2523), .B1(n792), .Y(n2524) );
  AOI22X1 U2223 ( .A0(n942), .A1(n886), .B0(n2809), .B1(n882), .Y(n2810) );
  AOI22X1 U2224 ( .A0(n1101), .A1(n1045), .B0(n3043), .B1(n1041), .Y(n3044) );
  AOI22X1 U2225 ( .A0(n624), .A1(n568), .B0(n3511), .B1(n564), .Y(n3512) );
  AOI22X1 U2226 ( .A0(n783), .A1(n727), .B0(n2575), .B1(n723), .Y(n2576) );
  XOR2X1 U2227 ( .A(n951), .B(n2757), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128224392_128224616_128224784)
         );
  XOR2X1 U2228 ( .A(n1110), .B(n2991), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128224392_128224616_128224784)
         );
  XOR2X1 U2229 ( .A(n633), .B(n3459), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128224392_128224616_128224784)
         );
  XOR2X1 U2230 ( .A(n792), .B(n2523), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128224392_128224616_128224784)
         );
  XOR2X1 U2231 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .Y(n2995) );
  XOR2X1 U2232 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .Y(n3463) );
  XOR2X1 U2233 ( .A(n904), .B(n932), .Y(n2751) );
  XOR2X1 U2234 ( .A(n1063), .B(n1091), .Y(n2985) );
  XOR2X1 U2235 ( .A(n586), .B(n614), .Y(n3453) );
  XOR2X1 U2236 ( .A(n745), .B(n773), .Y(n2517) );
  XOR2X1 U2237 ( .A(n902), .B(n923), .Y(n2757) );
  XOR2X1 U2238 ( .A(n1061), .B(n1082), .Y(n2991) );
  XOR2X1 U2239 ( .A(n584), .B(n605), .Y(n3459) );
  XOR2X1 U2240 ( .A(n743), .B(n764), .Y(n2523) );
  XOR2X1 U2241 ( .A(n886), .B(n942), .Y(n2809) );
  XOR2X1 U2242 ( .A(n1045), .B(n1101), .Y(n3043) );
  XOR2X1 U2243 ( .A(n568), .B(n624), .Y(n3511) );
  XOR2X1 U2244 ( .A(n727), .B(n783), .Y(n2575) );
  XOR2X1 U2245 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127827752_127827920)
         );
  XOR2X1 U2246 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127731920_127721600), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127672896_127674800_127730016), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127827752_127827920)
         );
  XOR2X1 U2247 ( .A(n962), .B(n2751), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128223720_128223944_128224168)
         );
  XOR2X1 U2248 ( .A(n1121), .B(n2985), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128223720_128223944_128224168)
         );
  XOR2X1 U2249 ( .A(n644), .B(n3453), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128223720_128223944_128224168)
         );
  XOR2X1 U2250 ( .A(n803), .B(n2517), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128223720_128223944_128224168)
         );
  XOR2X1 U2251 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128198024_128197968)
         );
  XOR2X1 U2252 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128198024_128197968)
         );
  XOR2X1 U2253 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128198024_128197968)
         );
  XOR2X1 U2254 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128198024_128197968) );
  XOR2X1 U2255 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .B(n2723), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127826576_127826800_127826968)
         );
  XOR2X1 U2256 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .B(n2957), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127826576_127826800_127826968)
         );
  XOR2X1 U2257 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .B(n3425), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127826576_127826800_127826968)
         );
  XOR2X1 U2258 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127830672_127844928_127846832), 
        .B(n2489), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127826576_127826800_127826968)
         );
  XOR2X1 U2259 ( .A(n976), .B(n2741), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128222376_128222600_128222768)
         );
  XOR2X1 U2260 ( .A(n1135), .B(n2975), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128222376_128222600_128222768)
         );
  XOR2X1 U2261 ( .A(n658), .B(n3443), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128222376_128222600_128222768)
         );
  XOR2X1 U2262 ( .A(n817), .B(n2507), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128222376_128222600_128222768)
         );
  XOR2X1 U2263 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .B(n2767), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128197520_128197632_128197800)
         );
  XOR2X1 U2264 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .B(n2533), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128197520_128197632_128197800)
         );
  XOR2X1 U2265 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .B(n2771), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128198080_128198192_128198360)
         );
  XOR2X1 U2266 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .B(n3005), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128198080_128198192_128198360)
         );
  XOR2X1 U2267 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .B(n3473), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128198080_128198192_128198360)
         );
  XOR2X1 U2268 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127831904_127846160_127848064), 
        .B(n2537), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128198080_128198192_128198360)
         );
  OR3XL U2269 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[3]), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[4]), .C(n3717), 
        .Y(n3715) );
  OR3XL U2270 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[3]), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[4]), .C(n3765), 
        .Y(n3763) );
  OR3XL U2271 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[3]), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[4]), .C(n3861), 
        .Y(n3859) );
  OR3XL U2272 ( .A(input_times_b0_mul_componentxUMxfirst_vector[3]), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[4]), .C(n3669), 
        .Y(n3667) );
  XOR2X1 U2273 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .B(n2773), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128198472_128198640_128198808)
         );
  XOR2X1 U2274 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .B(n3007), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128198472_128198640_128198808)
         );
  XOR2X1 U2275 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .B(n3475), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128198472_128198640_128198808)
         );
  XOR2X1 U2276 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .B(n2539), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128198472_128198640_128198808)
         );
  AND2X2 U2277 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer2_128198024_128197968)
         );
  AND2X2 U2278 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer2_128198024_128197968)
         );
  AND2X2 U2279 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer2_128198024_128197968)
         );
  AND2X2 U2280 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127715760_127848800_127850704), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127636256_127638160_127713856), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer2_128198024_128197968)
         );
  INVX1 U2281 ( .A(n4444), .Y(n957) );
  AOI22X1 U2282 ( .A0(n2311), .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[7]), 
        .B1(n4442), .Y(n4444) );
  XOR2X1 U2283 ( .A(n3713), .B(n2311), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[7]) );
  INVX1 U2284 ( .A(input_times_b0_mul_componentxn93), .Y(n798) );
  AOI22X1 U2285 ( .A0(input_times_b0_mul_componentxUMxAdder_finalxn47), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[7]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn93) );
  XOR2X1 U2286 ( .A(n3665), 
        .B(input_times_b0_mul_componentxUMxAdder_finalxn47), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[7]) );
  AND2X2 U2287 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer2_127826128_127826296)
         );
  AND2X2 U2288 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer2_127826128_127826296)
         );
  AND2X2 U2289 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer2_127826128_127826296)
         );
  AND2X2 U2290 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(input_times_b0_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer2_127826128_127826296)
         );
  AND2X2 U2291 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n987), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer3_128246112_128246336)
         );
  AND2X2 U2292 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n1146), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer3_128246112_128246336)
         );
  AND2X2 U2293 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n669), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer3_128246112_128246336)
         );
  AND2X2 U2294 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n828), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer3_128246112_128246336)
         );
  INVX1 U2295 ( .A(n4446), .Y(n972) );
  AOI22X1 U2296 ( .A0(input_p1_times_b1_mul_componentxUMxfirst_vector[5]), 
        .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[5]), 
        .B1(n4442), .Y(n4446) );
  XOR2X1 U2297 ( .A(n3715), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[5]), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[5]) );
  INVX1 U2298 ( .A(input_times_b0_mul_componentxn95), .Y(n813) );
  AOI22X1 U2299 ( .A0(input_times_b0_mul_componentxUMxfirst_vector[5]), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[5]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn95) );
  XOR2X1 U2300 ( .A(n3667), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[5]), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[5]) );
  INVX1 U2301 ( .A(n4443), .Y(n950) );
  AOI22X1 U2302 ( .A0(input_p1_times_b1_mul_componentxunsigned_output_8), 
        .A1(n125), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[8]), 
        .B1(n4442), .Y(n4443) );
  XOR2X1 U2303 ( .A(n3712), 
        .B(input_p1_times_b1_mul_componentxunsigned_output_8), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[8]) );
  OR2X2 U2304 ( .A(n2311), .B(n3713), .Y(n3712) );
  INVX1 U2305 ( .A(n4496), .Y(n1109) );
  AOI22X1 U2306 ( .A0(input_p2_times_b2_mul_componentxunsigned_output_8), 
        .A1(n129), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[8]), 
        .B1(n4495), .Y(n4496) );
  XOR2X1 U2307 ( .A(n3760), 
        .B(input_p2_times_b2_mul_componentxunsigned_output_8), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[8]) );
  OR2X2 U2308 ( .A(n2332), .B(n3761), .Y(n3760) );
  INVX1 U2309 ( .A(n4602), .Y(n632) );
  AOI22X1 U2310 ( .A0(output_p2_times_a2_mul_componentxunsigned_output_8), 
        .A1(n117), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[8]), 
        .B1(n4601), .Y(n4602) );
  XOR2X1 U2311 ( .A(n3856), 
        .B(output_p2_times_a2_mul_componentxunsigned_output_8), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[8]) );
  OR2X2 U2312 ( .A(n2374), .B(n3857), .Y(n3856) );
  INVX1 U2313 ( .A(input_times_b0_mul_componentxn92), .Y(n791) );
  AOI22X1 U2314 ( .A0(input_times_b0_mul_componentxunsigned_output_8), 
        .A1(n121), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[8]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn92) );
  XOR2X1 U2315 ( .A(n3664), .B(input_times_b0_mul_componentxunsigned_output_8), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[8]) );
  OR2X2 U2316 ( .A(input_times_b0_mul_componentxUMxAdder_finalxn47), .B(n3665), 
        .Y(n3664) );
  XOR2X1 U2317 ( 
        .A(input_p1_times_b1_mul_componentxUMxcarry_layer2_128198976_128199144), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer2_128198304_128198528_128198696), 
        .Y(n2814) );
  XOR2X1 U2318 ( .A(n922), .B(n2775), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128198304_128198528_128198696)
         );
  AND2X2 U2319 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer2_128198976_128199144)
         );
  XOR2X1 U2320 ( .A(n921), .B(n877), .Y(n2775) );
  XOR2X1 U2321 ( 
        .A(input_p2_times_b2_mul_componentxUMxcarry_layer2_128198976_128199144), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer2_128198304_128198528_128198696), 
        .Y(n3048) );
  XOR2X1 U2322 ( .A(n1081), .B(n3009), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128198304_128198528_128198696)
         );
  AND2X2 U2323 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer2_128198976_128199144)
         );
  XOR2X1 U2324 ( .A(n1080), .B(n1036), .Y(n3009) );
  XOR2X1 U2325 ( 
        .A(output_p2_times_a2_mul_componentxUMxcarry_layer2_128198976_128199144), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer2_128198304_128198528_128198696), 
        .Y(n3516) );
  XOR2X1 U2326 ( .A(n604), .B(n3477), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128198304_128198528_128198696)
         );
  AND2X2 U2327 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer2_128198976_128199144)
         );
  XOR2X1 U2328 ( .A(n603), .B(n559), .Y(n3477) );
  XOR2X1 U2329 ( 
        .A(input_times_b0_mul_componentxUMxcarry_layer2_128198976_128199144), 
        .B(input_times_b0_mul_componentxUMxsum_layer2_128198304_128198528_128198696), 
        .Y(n2580) );
  XOR2X1 U2330 ( .A(n763), .B(n2541), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128198304_128198528_128198696)
         );
  AND2X2 U2331 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer2_128198976_128199144)
         );
  XOR2X1 U2332 ( .A(n762), .B(n718), .Y(n2541) );
  XOR2X1 U2333 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128198976_128199144)
         );
  XOR2X1 U2334 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128198976_128199144)
         );
  XOR2X1 U2335 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128198976_128199144)
         );
  XOR2X1 U2336 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127627504_127629408), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127715872_127848912_127850816), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128198976_128199144) );
  XOR2X1 U2337 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127672560_127674464), 
        .B(n2721), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127826464_127826632_127826744)
         );
  XOR2X1 U2338 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .B(n2719), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_127672448_127826240_127826520)
         );
  XOR2X1 U2339 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127672560_127674464), 
        .B(n2955), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127826464_127826632_127826744)
         );
  XOR2X1 U2340 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .B(n2953), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_127672448_127826240_127826520)
         );
  XOR2X1 U2341 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127672560_127674464), 
        .B(n3423), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127826464_127826632_127826744)
         );
  XOR2X1 U2342 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .B(n3421), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_127672448_127826240_127826520)
         );
  XOR2X1 U2343 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127672560_127674464), 
        .B(n2487), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127826464_127826632_127826744)
         );
  XOR2X1 U2344 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .B(n2485), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_127672448_127826240_127826520)
         );
  XOR2X1 U2345 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n987), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer3_128246112_128246336)
         );
  XOR2X1 U2346 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n1146), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer3_128246112_128246336)
         );
  XOR2X1 U2347 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n669), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer3_128246112_128246336)
         );
  XOR2X1 U2348 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer2_127826464_127826632_127826744), 
        .B(n828), 
        .Y(input_times_b0_mul_componentxUMxsum_layer3_128246112_128246336) );
  INVX1 U2349 ( .A(n4445), .Y(n965) );
  AOI22X1 U2350 ( .A0(input_p1_times_b1_mul_componentxUMxfirst_vector[6]), 
        .A1(n125), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[6]), 
        .B1(n4442), .Y(n4445) );
  XOR2X1 U2351 ( .A(n3714), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[6]), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[6]) );
  OR2X2 U2352 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[5]), 
        .B(n3715), .Y(n3714) );
  INVX1 U2353 ( .A(n4498), .Y(n1124) );
  AOI22X1 U2354 ( .A0(input_p2_times_b2_mul_componentxUMxfirst_vector[6]), 
        .A1(n129), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[6]), 
        .B1(n4495), .Y(n4498) );
  XOR2X1 U2355 ( .A(n3762), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[6]), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[6]) );
  OR2X2 U2356 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[5]), 
        .B(n3763), .Y(n3762) );
  INVX1 U2357 ( .A(n4604), .Y(n647) );
  AOI22X1 U2358 ( .A0(output_p2_times_a2_mul_componentxUMxfirst_vector[6]), 
        .A1(n117), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[6]), 
        .B1(n4601), .Y(n4604) );
  XOR2X1 U2359 ( .A(n3858), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[6]), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[6]) );
  OR2X2 U2360 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[5]), 
        .B(n3859), .Y(n3858) );
  INVX1 U2361 ( .A(input_times_b0_mul_componentxn94), .Y(n806) );
  AOI22X1 U2362 ( .A0(input_times_b0_mul_componentxUMxfirst_vector[6]), 
        .A1(n121), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[6]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn94) );
  XOR2X1 U2363 ( .A(n3666), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[6]), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[6]) );
  OR2X2 U2364 ( .A(input_times_b0_mul_componentxUMxfirst_vector[5]), .B(n3667), 
        .Y(n3666) );
  INVX1 U2365 ( .A(n2752), .Y(n903) );
  AOI22X1 U2366 ( .A0(n932), .A1(n904), .B0(n2751), .B1(n962), .Y(n2752) );
  INVX1 U2367 ( .A(n2986), .Y(n1062) );
  AOI22X1 U2368 ( .A0(n1091), .A1(n1063), .B0(n2985), .B1(n1121), .Y(n2986) );
  INVX1 U2369 ( .A(n3454), .Y(n585) );
  AOI22X1 U2370 ( .A0(n614), .A1(n586), .B0(n3453), .B1(n644), .Y(n3454) );
  INVX1 U2371 ( .A(n2518), .Y(n744) );
  AOI22X1 U2372 ( .A0(n773), .A1(n745), .B0(n2517), .B1(n803), .Y(n2518) );
  INVX1 U2373 ( .A(n2766), .Y(n942) );
  AOI22X1 U2374 ( .A0(n967), .A1(n943), .B0(n2765), .B1(n991), .Y(n2766) );
  INVX1 U2375 ( .A(n3000), .Y(n1101) );
  AOI22X1 U2376 ( .A0(n1126), .A1(n1102), .B0(n2999), .B1(n1150), .Y(n3000) );
  INVX1 U2377 ( .A(n3468), .Y(n624) );
  AOI22X1 U2378 ( .A0(n649), .A1(n625), .B0(n3467), .B1(n673), .Y(n3468) );
  INVX1 U2379 ( .A(n2532), .Y(n783) );
  AOI22X1 U2380 ( .A0(n808), .A1(n784), .B0(n2531), .B1(n832), .Y(n2532) );
  INVX1 U2381 ( .A(n2762), .Y(n889) );
  AOI22X1 U2382 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B0(n2761), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .Y(n2762) );
  INVX1 U2383 ( .A(n2996), .Y(n1048) );
  AOI22X1 U2384 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B0(n2995), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .Y(n2996) );
  INVX1 U2385 ( .A(n3464), .Y(n571) );
  AOI22X1 U2386 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B0(n3463), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .Y(n3464) );
  INVX1 U2387 ( .A(n2528), .Y(n730) );
  AOI22X1 U2388 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127732704_127722384_127724288), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127673680_127675584_127730800), 
        .B0(n2527), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127636144_127638048_127713744), 
        .Y(n2528) );
  INVX1 U2389 ( .A(n2774), .Y(n874) );
  AOI22X1 U2390 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B0(n2773), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .Y(n2774) );
  INVX1 U2391 ( .A(n2540), .Y(n715) );
  AOI22X1 U2392 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B0(n2539), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127636368_127638272_127713968), 
        .Y(n2540) );
  XOR2X1 U2393 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(input_p1_times_b1_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[2]) );
  XOR2X1 U2394 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(input_p2_times_b2_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[2]) );
  XOR2X1 U2395 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(output_p2_times_a2_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[2]) );
  XOR2X1 U2396 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127830336_127844592_127846496), 
        .B(input_times_b0_mul_componentxUMxcarry_layer1_127830168_127844480), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[2]) );
  XOR2X1 U2397 ( .A(n931), .B(n2769), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128197464_128197688_128197856)
         );
  XOR2X1 U2398 ( .A(n1090), .B(n3003), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128197464_128197688_128197856)
         );
  XOR2X1 U2399 ( .A(n613), .B(n3471), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128197464_128197688_128197856)
         );
  XOR2X1 U2400 ( .A(n772), .B(n2535), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128197464_128197688_128197856)
         );
  XOR2X1 U2401 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .Y(n2767) );
  XOR2X1 U2402 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .Y(n3001) );
  XOR2X1 U2403 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .Y(n3469) );
  XOR2X1 U2404 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .Y(n2533) );
  XOR2X1 U2405 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .Y(n2773) );
  XOR2X1 U2406 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .Y(n3007) );
  XOR2X1 U2407 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .Y(n3475) );
  XOR2X1 U2408 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127673904_127675808_127731024), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127732928_127722608_127724512), 
        .Y(n2539) );
  XOR2X1 U2409 ( .A(n920), .B(n879), .Y(n2769) );
  XOR2X1 U2410 ( .A(n1079), .B(n1038), .Y(n3003) );
  XOR2X1 U2411 ( .A(n602), .B(n561), .Y(n3471) );
  XOR2X1 U2412 ( .A(n761), .B(n720), .Y(n2535) );
  XOR2X1 U2413 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .B(n3001), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128197520_128197632_128197800)
         );
  XOR2X1 U2414 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .B(n3469), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128197520_128197632_128197800)
         );
  OR3XL U2415 ( .A(n994), .B(n993), .C(n995), .Y(n3917) );
  OR3XL U2416 ( .A(n1153), .B(n1152), .C(n1154), .Y(n3960) );
  OR3XL U2417 ( .A(n676), .B(n675), .C(n677), .Y(n4046) );
  OR3XL U2418 ( .A(n835), .B(n834), .C(n836), .Y(n3874) );
  INVX1 U2419 ( .A(n4448), .Y(n986) );
  AOI22XL U2420 ( .A0(input_p1_times_b1_mul_componentxUMxfirst_vector[3]), 
        .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[3]), 
        .B1(n4442), .Y(n4448) );
  XOR2X1 U2421 ( .A(n3717), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[3]), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[3]) );
  INVX1 U2422 ( .A(n4501), .Y(n1145) );
  AOI22X1 U2423 ( .A0(input_p2_times_b2_mul_componentxUMxfirst_vector[3]), 
        .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[3]), 
        .B1(n4495), .Y(n4501) );
  XOR2X1 U2424 ( .A(n3765), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[3]), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[3]) );
  INVX1 U2425 ( .A(n4499), .Y(n1131) );
  AOI22XL U2426 ( .A0(input_p2_times_b2_mul_componentxUMxfirst_vector[5]), 
        .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[5]), 
        .B1(n4495), .Y(n4499) );
  XOR2X1 U2427 ( .A(n3763), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[5]), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[5]) );
  INVX1 U2428 ( .A(n4607), .Y(n668) );
  AOI22X1 U2429 ( .A0(output_p2_times_a2_mul_componentxUMxfirst_vector[3]), 
        .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[3]), 
        .B1(n4601), .Y(n4607) );
  XOR2X1 U2430 ( .A(n3861), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[3]), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[3]) );
  INVX1 U2431 ( .A(n4605), .Y(n654) );
  AOI22XL U2432 ( .A0(output_p2_times_a2_mul_componentxUMxfirst_vector[5]), 
        .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[5]), 
        .B1(n4601), .Y(n4605) );
  XOR2X1 U2433 ( .A(n3859), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[5]), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[5]) );
  INVX1 U2434 ( .A(input_times_b0_mul_componentxn97), .Y(n827) );
  AOI22XL U2435 ( .A0(input_times_b0_mul_componentxUMxfirst_vector[3]), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[3]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn97) );
  XOR2X1 U2436 ( .A(n3669), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[3]), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[3]) );
  INVX1 U2437 ( .A(n4447), .Y(n980) );
  AOI22XL U2438 ( .A0(input_p1_times_b1_mul_componentxUMxfirst_vector[4]), 
        .A1(n125), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[4]), 
        .B1(n4442), .Y(n4447) );
  XOR2X1 U2439 ( .A(n3716), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[4]), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[4]) );
  OR2X2 U2440 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[3]), 
        .B(n3717), .Y(n3716) );
  INVX1 U2441 ( .A(n4500), .Y(n1139) );
  AOI22XL U2442 ( .A0(input_p2_times_b2_mul_componentxUMxfirst_vector[4]), 
        .A1(n129), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[4]), 
        .B1(n4495), .Y(n4500) );
  XOR2X1 U2443 ( .A(n3764), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[4]), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[4]) );
  OR2X2 U2444 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[3]), 
        .B(n3765), .Y(n3764) );
  INVX1 U2445 ( .A(n4606), .Y(n662) );
  AOI22XL U2446 ( .A0(output_p2_times_a2_mul_componentxUMxfirst_vector[4]), 
        .A1(n117), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[4]), 
        .B1(n4601), .Y(n4606) );
  XOR2X1 U2447 ( .A(n3860), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[4]), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[4]) );
  OR2X2 U2448 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[3]), 
        .B(n3861), .Y(n3860) );
  INVX1 U2449 ( .A(input_times_b0_mul_componentxn96), .Y(n821) );
  AOI22XL U2450 ( .A0(input_times_b0_mul_componentxUMxfirst_vector[4]), 
        .A1(n121), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[4]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn96) );
  XOR2X1 U2451 ( .A(n3668), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[4]), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[4]) );
  OR2X2 U2452 ( .A(input_times_b0_mul_componentxUMxfirst_vector[3]), .B(n3669), 
        .Y(n3668) );
  INVX1 U2453 ( .A(n2768), .Y(n882) );
  AOI22X1 U2454 ( 
        .A0(input_p1_times_b1_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .A1(input_p1_times_b1_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B0(n2767), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .Y(n2768) );
  INVX1 U2455 ( .A(n3002), .Y(n1041) );
  AOI22X1 U2456 ( 
        .A0(input_p2_times_b2_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .A1(input_p2_times_b2_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B0(n3001), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .Y(n3002) );
  INVX1 U2457 ( .A(n3470), .Y(n564) );
  AOI22X1 U2458 ( 
        .A0(output_p2_times_a2_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .A1(output_p2_times_a2_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B0(n3469), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .Y(n3470) );
  INVX1 U2459 ( .A(n2534), .Y(n723) );
  AOI22X1 U2460 ( 
        .A0(input_times_b0_mul_componentxUMxsum_layer1_127673792_127675696_127730912), 
        .A1(input_times_b0_mul_componentxUMxsum_layer1_127831792_127846048_127847952), 
        .B0(n2533), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127732816_127722496_127724400), 
        .Y(n2534) );
  XNOR2X1 U2461 ( .A(n993), .B(n3918), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[2]) );
  NOR2X1 U2462 ( .A(n995), .B(n994), .Y(n3918) );
  XNOR2X1 U2463 ( .A(n1152), .B(n3961), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[2]) );
  NOR2X1 U2464 ( .A(n1154), .B(n1153), .Y(n3961) );
  XNOR2X1 U2465 ( .A(n675), .B(n4047), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[2]) );
  NOR2X1 U2466 ( .A(n677), .B(n676), .Y(n4047) );
  XNOR2X1 U2467 ( .A(n834), .B(n3875), 
        .Y(input_times_b0_div_componentxinput_A_inverted[2]) );
  NOR2X1 U2468 ( .A(n836), .B(n835), .Y(n3875) );
  XOR2X1 U2469 ( .A(n994), .B(n995), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[1]) );
  XOR2X1 U2470 ( .A(n1153), .B(n1154), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[1]) );
  XOR2X1 U2471 ( .A(n676), .B(n677), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[1]) );
  XOR2X1 U2472 ( .A(n835), .B(n836), 
        .Y(input_times_b0_div_componentxinput_A_inverted[1]) );
  INVX1 U2473 ( .A(n258), .Y(n320) );
  INVX1 U2474 ( .A(n258), .Y(n319) );
  INVX1 U2475 ( .A(n258), .Y(n321) );
  BUFX3 U2476 ( .A(n161), .Y(n159) );
  BUFX3 U2477 ( .A(n161), .Y(n160) );
  BUFX3 U2478 ( .A(n162), .Y(n157) );
  BUFX3 U2479 ( .A(n162), .Y(n158) );
  BUFX3 U2480 ( .A(n163), .Y(n155) );
  BUFX3 U2481 ( .A(n163), .Y(n156) );
  BUFX3 U2482 ( .A(n164), .Y(n153) );
  BUFX3 U2483 ( .A(n164), .Y(n154) );
  BUFX3 U2484 ( .A(n257), .Y(n137) );
  BUFX3 U2485 ( .A(n257), .Y(n138) );
  NOR3X1 U2486 ( .A(n853), .B(n854), 
        .C(input_times_b0_div_componentxUDxinverter_for_substractionxn4), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn2) );
  NOR3X1 U2487 ( .A(n1012), .B(n1013), .C(n1762), .Y(n1761) );
  NOR3X1 U2488 ( .A(n1171), .B(n1172), .C(n1771), .Y(n1770) );
  NOR3X1 U2489 ( .A(n535), .B(n536), .C(n1780), .Y(n1779) );
  NOR3X1 U2490 ( .A(n694), .B(n695), .C(n1789), .Y(n1788) );
  NOR3X1 U2491 ( .A(output_contracterxn7), .B(output_previous_1[16]), 
        .C(output_previous_1[15]), .Y(output_contracterxn2) );
  OR3XL U2492 ( .A(n165), .B(output_previous_1[8]), .C(output_previous_1[9]), 
        .Y(output_contracterxn7) );
  XOR2X1 U2493 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn16), 
        .B(n838), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[11]) );
  XOR2X1 U2494 ( .A(n1768), .B(n997), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[11])
         );
  XOR2X1 U2495 ( .A(n1777), .B(n1156), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[11])
         );
  XOR2X1 U2496 ( .A(n1786), .B(n520), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[11])
         );
  XOR2X1 U2497 ( .A(n1795), .B(n679), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[11])
         );
  XOR2X1 U2498 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn4), 
        .B(n853), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[7]) );
  XOR2X1 U2499 ( .A(n1762), .B(n1012), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[7])
         );
  XOR2X1 U2500 ( .A(n1771), .B(n1171), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[7])
         );
  XOR2X1 U2501 ( .A(n1780), .B(n535), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[7])
         );
  XOR2X1 U2502 ( .A(n1789), .B(n694), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[7])
         );
  XOR2X1 U2503 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn14), 
        .B(n840), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[13]) );
  XOR2X1 U2504 ( .A(n1767), .B(n999), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[13])
         );
  XOR2X1 U2505 ( .A(n1776), .B(n1158), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[13])
         );
  XOR2X1 U2506 ( .A(n1785), .B(n522), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[13])
         );
  XOR2X1 U2507 ( .A(n1794), .B(n681), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[13])
         );
  XOR2X1 U2508 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn12), 
        .B(n842), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[15]) );
  XOR2X1 U2509 ( .A(n1766), .B(n1001), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[15])
         );
  XOR2X1 U2510 ( .A(n1775), .B(n1160), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[15])
         );
  XOR2X1 U2511 ( .A(n1784), .B(n524), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[15])
         );
  XOR2X1 U2512 ( .A(n1793), .B(n683), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[15])
         );
  XNOR2X1 U2513 ( .A(n64), .B(n854), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[8]) );
  NOR2X1 U2514 ( .A(n853), 
        .B(input_times_b0_div_componentxUDxinverter_for_substractionxn4), 
        .Y(n64) );
  XNOR2X1 U2515 ( .A(n65), .B(n1013), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[8])
         );
  NOR2X1 U2516 ( .A(n1012), .B(n1762), .Y(n65) );
  XNOR2X1 U2517 ( .A(n66), .B(n1172), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[8])
         );
  NOR2X1 U2518 ( .A(n1171), .B(n1771), .Y(n66) );
  XNOR2X1 U2519 ( .A(n67), .B(n536), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[8])
         );
  NOR2X1 U2520 ( .A(n535), .B(n1780), .Y(n67) );
  XNOR2X1 U2521 ( .A(n68), .B(n695), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[8])
         );
  NOR2X1 U2522 ( .A(n694), .B(n1789), .Y(n68) );
  XNOR2X1 U2523 ( .A(n69), .B(n839), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[12]) );
  NOR2X1 U2524 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn16), 
        .B(n838), .Y(n69) );
  XNOR2X1 U2525 ( .A(n70), .B(n998), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[12])
         );
  NOR2X1 U2526 ( .A(n1768), .B(n997), .Y(n70) );
  XNOR2X1 U2527 ( .A(n71), .B(n1157), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[12])
         );
  NOR2X1 U2528 ( .A(n1777), .B(n1156), .Y(n71) );
  XNOR2X1 U2529 ( .A(n72), .B(n521), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[12])
         );
  NOR2X1 U2530 ( .A(n1786), .B(n520), .Y(n72) );
  XNOR2X1 U2531 ( .A(n73), .B(n680), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[12])
         );
  NOR2X1 U2532 ( .A(n1795), .B(n679), .Y(n73) );
  XNOR2X1 U2533 ( .A(n74), .B(n841), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[14]) );
  NOR2X1 U2534 ( .A(n840), 
        .B(input_times_b0_div_componentxUDxinverter_for_substractionxn14), 
        .Y(n74) );
  XNOR2X1 U2535 ( .A(n75), .B(n1000), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[14])
         );
  NOR2X1 U2536 ( .A(n999), .B(n1767), .Y(n75) );
  XNOR2X1 U2537 ( .A(n76), .B(n1159), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[14])
         );
  NOR2X1 U2538 ( .A(n1158), .B(n1776), .Y(n76) );
  XNOR2X1 U2539 ( .A(n77), .B(n523), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[14])
         );
  NOR2X1 U2540 ( .A(n522), .B(n1785), .Y(n77) );
  XNOR2X1 U2541 ( .A(n78), .B(n682), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[14])
         );
  NOR2X1 U2542 ( .A(n681), .B(n1794), .Y(n78) );
  OR3XL U2543 ( .A(n838), .B(n839), 
        .C(input_times_b0_div_componentxUDxinverter_for_substractionxn16), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn14) );
  OR3XL U2544 ( .A(n997), .B(n998), .C(n1768), .Y(n1767) );
  OR3XL U2545 ( .A(n1156), .B(n1157), .C(n1777), .Y(n1776) );
  OR3XL U2546 ( .A(n520), .B(n521), .C(n1786), .Y(n1785) );
  OR3XL U2547 ( .A(n679), .B(n680), .C(n1795), .Y(n1794) );
  NAND3X1 U2548 ( .A(output_previous_1[16]), .B(output_previous_1[15]), 
        .C(n165), .Y(output_contracterxn6) );
  OR3XL U2549 ( .A(n840), .B(n841), 
        .C(input_times_b0_div_componentxUDxinverter_for_substractionxn14), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn12) );
  OR3XL U2550 ( .A(n999), .B(n1000), .C(n1767), .Y(n1766) );
  OR3XL U2551 ( .A(n1158), .B(n1159), .C(n1776), .Y(n1775) );
  OR3XL U2552 ( .A(n522), .B(n523), .C(n1785), .Y(n1784) );
  OR3XL U2553 ( .A(n681), .B(n682), .C(n1794), .Y(n1793) );
  BUFX3 U2554 ( .A(output_previous_1[17]), .Y(n165) );
  XOR2X1 U2555 ( .A(n4169), .B(n4170), .Y(output_previous_1[17]) );
  XNOR2X1 U2556 ( .A(results_a1_a2_inv[17]), .B(results_b0_b1_b2[17]), 
        .Y(n4169) );
  AOI22X1 U2557 ( .A0(n4171), .A1(n1205), .B0(results_b0_b1_b2[16]), 
        .B1(results_a1_a2_inv[16]), .Y(n4170) );
  XOR2X1 U2558 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b4), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b3), .Y(n3095) );
  XOR2X1 U2559 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b5), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b4), .Y(n3097) );
  XOR2X1 U2560 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b0), .B(n494), 
        .Y(n3193) );
  XOR2X1 U2561 ( .A(n4121), .B(n4122), .Y(results_a1_a2[8]) );
  XOR2X1 U2562 ( .A(results_b0_b1_adderxn14), .B(results_b0_b1_adderxn15), 
        .Y(results_b0_b1[3]) );
  XOR2X1 U2563 ( .A(n4098), .B(n4099), .Y(results_b0_b1_b2[3]) );
  XOR2X1 U2564 ( .A(results_b0_b1_adderxn10), .B(results_b0_b1_adderxn11), 
        .Y(results_b0_b1[5]) );
  XOR2X1 U2565 ( .A(n4094), .B(n4095), .Y(results_b0_b1_b2[5]) );
  XOR2X1 U2566 ( .A(results_b0_b1_adderxn6), .B(results_b0_b1_adderxn7), 
        .Y(results_b0_b1[7]) );
  XOR2X1 U2567 ( .A(n4090), .B(n4091), .Y(results_b0_b1_b2[7]) );
  XOR2X1 U2568 ( .A(results_b0_b1_adderxn2), .B(results_b0_b1_adderxn3), 
        .Y(results_b0_b1[9]) );
  XOR2X1 U2569 ( .A(n4086), .B(n4087), .Y(results_b0_b1_b2[9]) );
  XOR2X1 U2570 ( .A(results_b0_b1_adderxn32), .B(results_b0_b1_adderxn33), 
        .Y(results_b0_b1[11]) );
  XOR2X1 U2571 ( .A(n4115), .B(n4116), .Y(results_b0_b1_b2[11]) );
  XOR2X1 U2572 ( .A(results_b0_b1_adderxn28), .B(results_b0_b1_adderxn29), 
        .Y(results_b0_b1[13]) );
  XOR2X1 U2573 ( .A(n4111), .B(n4112), .Y(results_b0_b1_b2[13]) );
  XOR2X1 U2574 ( .A(n4107), .B(n4108), .Y(results_b0_b1_b2[15]) );
  XOR2X1 U2575 ( .A(n4125), .B(n4126), .Y(results_a1_a2[6]) );
  XOR2X1 U2576 ( .A(results_b0_b1_adderxn16), .B(results_b0_b1_adderxn17), 
        .Y(results_b0_b1[2]) );
  XOR2X1 U2577 ( .A(n4100), .B(n4101), .Y(results_b0_b1_b2[2]) );
  XOR2X1 U2578 ( .A(results_b0_b1_adderxn12), .B(results_b0_b1_adderxn13), 
        .Y(results_b0_b1[4]) );
  XOR2X1 U2579 ( .A(n4096), .B(n4097), .Y(results_b0_b1_b2[4]) );
  XOR2X1 U2580 ( .A(results_b0_b1_adderxn8), .B(results_b0_b1_adderxn9), 
        .Y(results_b0_b1[6]) );
  XOR2X1 U2581 ( .A(n4092), .B(n4093), .Y(results_b0_b1_b2[6]) );
  XOR2X1 U2582 ( .A(results_b0_b1_adderxn4), .B(results_b0_b1_adderxn5), 
        .Y(results_b0_b1[8]) );
  XOR2X1 U2583 ( .A(n4088), .B(n4089), .Y(results_b0_b1_b2[8]) );
  XOR2X1 U2584 ( .A(results_b0_b1_adderxn35), .B(results_b0_b1_adderxn34), 
        .Y(results_b0_b1[10]) );
  XOR2X1 U2585 ( .A(n4118), .B(n4117), .Y(results_b0_b1_b2[10]) );
  XOR2X1 U2586 ( .A(results_b0_b1_adderxn31), .B(results_b0_b1_adderxn30), 
        .Y(results_b0_b1[12]) );
  XOR2X1 U2587 ( .A(n4114), .B(n4113), .Y(results_b0_b1_b2[12]) );
  XOR2X1 U2588 ( .A(results_b0_b1_adderxn27), .B(results_b0_b1_adderxn26), 
        .Y(results_b0_b1[14]) );
  XOR2X1 U2589 ( .A(n4110), .B(n4109), .Y(results_b0_b1_b2[14]) );
  INVX1 U2590 ( .A(n3098), .Y(n494) );
  AOI22X1 U2591 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b4), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b5), .B0(n3097), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b3), .Y(n3098) );
  INVX1 U2592 ( .A(n3096), .Y(n501) );
  AOI22X1 U2593 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b3), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b4), .B0(n3095), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b2), .Y(n3096) );
  INVX1 U2594 ( .A(n3194), .Y(n493) );
  AOI22X1 U2595 ( .A0(n494), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b0), .B0(n3193), 
        .B1(n513), .Y(n3194) );
  BUFX3 U2596 ( .A(n1321), .Y(n146) );
  BUFX3 U2597 ( .A(n1341), .Y(n148) );
  BUFX3 U2598 ( .A(n1380), .Y(n152) );
  BUFX3 U2599 ( .A(n1238), .Y(n136) );
  AOI32X1 U2600 ( .A0(results_a1_a2_inv[0]), .A1(n4168), 
        .A2(results_b0_b1_b2[0]), .B0(results_a1_a2_inv[1]), 
        .B1(results_b0_b1_b2[1]), .Y(n4167) );
  NOR2X1 U2601 ( .A(n4528), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b10) );
  NOR2X1 U2602 ( .A(n4527), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b11) );
  NOR2X1 U2603 ( .A(n4526), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b12) );
  NOR2X1 U2604 ( .A(n214), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b7) );
  NOR2X1 U2605 ( .A(n213), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b8) );
  NOR2X1 U2606 ( .A(n212), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b9) );
  NOR2X1 U2607 ( .A(n213), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b8) );
  NOR2X1 U2608 ( .A(n214), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b7) );
  INVX1 U2609 ( .A(n3142), .Y(n504) );
  AOI22X1 U2610 ( .A0(output_p1_times_a1_mul_componentxUMxa10_and_b2), 
        .A1(output_p1_times_a1_mul_componentxUMxa9_and_b3), .B0(n3141), 
        .B1(output_p1_times_a1_mul_componentxUMxa11_and_b1), .Y(n3142) );
  NOR2X1 U2611 ( .A(n231), .B(n4528), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b10) );
  NOR2X1 U2612 ( .A(n231), .B(n4527), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b11) );
  INVX1 U2613 ( .A(n3094), .Y(n508) );
  AOI22X1 U2614 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b2), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b3), .B0(n3093), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b1), .Y(n3094) );
  INVX1 U2615 ( .A(n3108), .Y(n500) );
  AOI22X1 U2616 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b3), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b4), .B0(n3107), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b2), .Y(n3108) );
  INVX1 U2617 ( .A(n3106), .Y(n479) );
  AOI22X1 U2618 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b6), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b7), .B0(n3105), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b5), .Y(n3106) );
  INVX1 U2619 ( .A(n3092), .Y(n515) );
  AOI22X1 U2620 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b1), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b2), .B0(n3091), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b0), .Y(n3092) );
  INVX1 U2621 ( .A(n3102), .Y(n487) );
  AOI22X1 U2622 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b5), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b6), .B0(n3101), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b4), .Y(n3102) );
  INVX1 U2623 ( .A(n3110), .Y(n469) );
  AOI22X1 U2624 ( .A0(output_p1_times_a1_mul_componentxUMxa1_and_b7), 
        .A1(output_p1_times_a1_mul_componentxUMxa0_and_b8), .B0(n3109), 
        .B1(output_p1_times_a1_mul_componentxUMxa2_and_b6), .Y(n3110) );
  INVX1 U2625 ( .A(n3114), .Y(n512) );
  AOI22X1 U2626 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b1), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b2), .B0(n3113), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b0), .Y(n3114) );
  INVX1 U2627 ( .A(n3132), .Y(n491) );
  AOI22X1 U2628 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b4), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b5), .B0(n3131), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b3), .Y(n3132) );
  NOR2X1 U2629 ( .A(n231), .B(n4526), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b12) );
  NOR2X1 U2630 ( .A(n231), .B(n4525), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b13) );
  NOR2X1 U2631 ( .A(n231), .B(n214), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b7) );
  NOR2X1 U2632 ( .A(n231), .B(n213), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b8) );
  NOR2X1 U2633 ( .A(n231), .B(n212), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b9) );
  NOR2X1 U2634 ( .A(n212), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b9) );
  NOR2X1 U2635 ( .A(n214), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b7) );
  NOR2X1 U2636 ( .A(n214), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b7) );
  NOR2X1 U2637 ( .A(n213), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b8) );
  XOR2X1 U2638 ( .A(n4123), .B(n4124), .Y(results_a1_a2[7]) );
  XOR2X1 U2639 ( .A(n4144), .B(n4145), .Y(results_a1_a2[13]) );
  XOR2X1 U2640 ( .A(n4119), .B(n4120), .Y(results_a1_a2[9]) );
  XOR2X1 U2641 ( .A(n4131), .B(n4132), .Y(results_a1_a2[3]) );
  XOR2X1 U2642 ( .A(n4127), .B(n4128), .Y(results_a1_a2[5]) );
  XOR2X1 U2643 ( .A(n4148), .B(n4149), .Y(results_a1_a2[11]) );
  XOR2X1 U2644 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b2), .B(n3095), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127830560_127844816_127846720)
         );
  XOR2X1 U2645 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b3), .B(n3111), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673008_127674912_127730128)
         );
  XOR2X1 U2646 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b4), .B(n3139), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732480_127722160_127724064)
         );
  XOR2X1 U2647 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b5), .B(n3123), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673232_127675136_127730352)
         );
  XOR2X1 U2648 ( .A(output_p1_times_a1_mul_componentxUMxa12_and_b0), .B(n436), 
        .Y(n3213) );
  XOR2X1 U2649 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b3), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b2), .Y(n3093) );
  XOR2X1 U2650 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b7), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b6), .Y(n3105) );
  XOR2X1 U2651 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b2), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b1), .Y(n3091) );
  XOR2X1 U2652 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b6), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b5), .Y(n3101) );
  XOR2X1 U2653 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b0), .B(n515), 
        .Y(n3187) );
  XOR2X1 U2654 ( .A(output_p1_times_a1_mul_componentxUMxa9_and_b0), .B(n469), 
        .Y(n3201) );
  XOR2X1 U2655 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b2), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b1), .Y(n3099) );
  XOR2X1 U2656 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b2), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b1), .Y(n3113) );
  XOR2X1 U2657 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b3), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b2), .Y(n3103) );
  XOR2X1 U2658 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b3), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b2), .Y(n3119) );
  XOR2X1 U2659 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b4), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b3), .Y(n3107) );
  XOR2X1 U2660 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b4), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b3), .Y(n3125) );
  XOR2X1 U2661 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b5), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b4), .Y(n3111) );
  XOR2X1 U2662 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b5), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b4), .Y(n3131) );
  XOR2X1 U2663 ( .A(output_p1_times_a1_mul_componentxUMxa9_and_b2), 
        .B(output_p1_times_a1_mul_componentxUMxa10_and_b1), .Y(n3133) );
  XOR2X1 U2664 ( .A(output_p1_times_a1_mul_componentxUMxa9_and_b3), 
        .B(output_p1_times_a1_mul_componentxUMxa10_and_b2), .Y(n3141) );
  XOR2X1 U2665 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b6), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b5), .Y(n3117) );
  XOR2X1 U2666 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b7), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b6), .Y(n3123) );
  XOR2X1 U2667 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b6), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b5), .Y(n3139) );
  XOR2X1 U2668 ( .A(n4140), .B(n4141), .Y(results_a1_a2[15]) );
  XOR2X1 U2669 ( .A(n4143), .B(n4142), .Y(results_a1_a2[14]) );
  AND2X2 U2670 ( .A(output_p1_times_a1_mul_componentxUMxa4_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa3_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer1_127672560_127674464)
         );
  XOR2X1 U2671 ( .A(results_b0_b1_b2[1]), .B(results_a1_a2_inv[1]), .Y(n4168)
         );
  XOR2X1 U2672 ( .A(results_a1_a2[1]), .B(results_a1_a2_inv[0]), 
        .Y(results_a1_a2_inv[1]) );
  XNOR2X1 U2673 ( .A(results_a1_a2[2]), .B(results_a1_a2_inv_inverterxn9), 
        .Y(results_a1_a2_inv[2]) );
  NOR2X1 U2674 ( .A(results_a1_a2_inv[0]), .B(results_a1_a2[1]), 
        .Y(results_a1_a2_inv_inverterxn9) );
  XOR2X1 U2675 ( .A(results_b0_b1_adderxn24), .B(results_b0_b1_adderxn25), 
        .Y(results_b0_b1[15]) );
  XOR2X1 U2676 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b0), .B(n3099), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127672672_127674576_127729792)
         );
  XOR2X1 U2677 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b1), .B(n3119), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732144_127721824_127723728)
         );
  XOR2X1 U2678 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b6), .B(n3109), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127831008_127845264_127847168)
         );
  OR3XL U2679 ( .A(results_a1_a2[1]), .B(results_a1_a2[2]), 
        .C(results_a1_a2_inv[0]), .Y(results_a1_a2_inv_inverterxn8) );
  XOR2X1 U2680 ( .A(n4129), .B(n4130), .Y(results_a1_a2[4]) );
  XOR2X1 U2681 ( .A(n4147), .B(n4146), .Y(results_a1_a2[12]) );
  XOR2X1 U2682 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b0), .B(n3113), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732032_127721712_127723616)
         );
  XOR2X1 U2683 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b2), .B(n3125), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732256_127721936_127723840)
         );
  XOR2X1 U2684 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b3), .B(n3097), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127830672_127844928_127846832)
         );
  XOR2X1 U2685 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b4), .B(n3117), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673120_127675024_127730240)
         );
  XOR2X1 U2686 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b5), .B(n3105), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127830896_127845152_127847056)
         );
  XOR2X1 U2687 ( .A(output_p1_times_a1_mul_componentxUMxa4_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa3_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127672560_127674464)
         );
  XOR2X1 U2688 ( .A(results_b0_b1_adderxn22), .B(n1209), .Y(results_b0_b1[16])
         );
  XOR2X1 U2689 ( .A(n4105), .B(n1207), .Y(results_b0_b1_b2[16]) );
  XOR2X1 U2690 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b2), .B(n3107), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127672896_127674800_127730016)
         );
  XOR2X1 U2691 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b4), .B(n3101), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127830784_127845040_127846944)
         );
  XOR2X1 U2692 ( .A(n4151), .B(n4150), .Y(results_a1_a2[10]) );
  XOR2X1 U2693 ( .A(n4138), .B(n1301), .Y(results_a1_a2[16]) );
  AND2X2 U2694 ( .A(output_p1_times_a1_mul_componentxUMxa7_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa6_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer1_127731920_127721600)
         );
  XOR2X1 U2695 ( .A(n4133), .B(n4134), .Y(results_a1_a2[2]) );
  XOR2X1 U2696 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b1), .B(n3103), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127672784_127674688_127729904)
         );
  XOR2X1 U2697 ( .A(output_p1_times_a1_mul_componentxUMxa7_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa6_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127731920_127721600)
         );
  INVX1 U2698 ( .A(n3134), .Y(n511) );
  AOI22X1 U2699 ( .A0(output_p1_times_a1_mul_componentxUMxa10_and_b1), 
        .A1(output_p1_times_a1_mul_componentxUMxa9_and_b2), .B0(n3133), 
        .B1(output_p1_times_a1_mul_componentxUMxa11_and_b0), .Y(n3134) );
  INVX1 U2700 ( .A(n3104), .Y(n506) );
  AOI22X1 U2701 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b2), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b3), .B0(n3103), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b1), .Y(n3104) );
  INVX1 U2702 ( .A(n3118), .Y(n486) );
  AOI22X1 U2703 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b5), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b6), .B0(n3117), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b4), .Y(n3118) );
  INVX1 U2704 ( .A(n3202), .Y(n468) );
  AOI22X1 U2705 ( .A0(n469), 
        .A1(output_p1_times_a1_mul_componentxUMxa9_and_b0), .B0(n3201), 
        .B1(n492), .Y(n3202) );
  INVX1 U2706 ( .A(n3124), .Y(n476) );
  AOI22X1 U2707 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b6), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b7), .B0(n3123), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b5), .Y(n3124) );
  BUFX3 U2708 ( .A(n1321), .Y(n145) );
  BUFX3 U2709 ( .A(n1341), .Y(n147) );
  BUFX3 U2710 ( .A(n1380), .Y(n151) );
  BUFX3 U2711 ( .A(n1238), .Y(n135) );
  BUFX3 U2712 ( .A(n1360), .Y(n149) );
  INVX1 U2713 ( .A(n3214), .Y(n435) );
  AOI22X1 U2714 ( .A0(n436), 
        .A1(output_p1_times_a1_mul_componentxUMxa12_and_b0), .B0(n3213), 
        .B1(n467), .Y(n3214) );
  INVX1 U2715 ( .A(n3100), .Y(n513) );
  AOI22X1 U2716 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b1), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b2), .B0(n3099), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b0), .Y(n3100) );
  INVX1 U2717 ( .A(n3112), .Y(n492) );
  AOI22X1 U2718 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b4), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b5), .B0(n3111), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b3), .Y(n3112) );
  INVX1 U2719 ( .A(n3130), .Y(n467) );
  AOI22X1 U2720 ( .A0(output_p1_times_a1_mul_componentxUMxa4_and_b7), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b8), .B0(n3129), 
        .B1(output_p1_times_a1_mul_componentxUMxa5_and_b6), .Y(n3130) );
  INVX1 U2721 ( .A(n3120), .Y(n505) );
  AOI22X1 U2722 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b2), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b3), .B0(n3119), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b1), .Y(n3120) );
  INVX1 U2723 ( .A(n3188), .Y(n510) );
  AOI22X1 U2724 ( .A0(n515), 
        .A1(output_p1_times_a1_mul_componentxUMxa3_and_b0), .B0(n3187), 
        .B1(output_p1_times_a1_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .Y(n3188) );
  BUFX3 U2725 ( .A(n1360), .Y(n150) );
  NAND2X1 U2726 ( .A(results_b0_b1_b2[0]), .B(results_a1_a2_inv[0]), .Y(n79)
         );
  NOR2X1 U2727 ( .A(n4528), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b10) );
  NOR2X1 U2728 ( .A(n4527), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b11) );
  NOR2X1 U2729 ( .A(n4525), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b13) );
  NOR2X1 U2730 ( .A(n4524), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b14) );
  NOR2X1 U2731 ( .A(n212), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b9) );
  NOR2X1 U2732 ( .A(n214), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b7) );
  NOR2X1 U2733 ( .A(n4528), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b10) );
  INVX1 U2734 ( .A(n3150), .Y(n498) );
  AOI22X1 U2735 ( .A0(output_p1_times_a1_mul_componentxUMxa10_and_b3), 
        .A1(output_p1_times_a1_mul_componentxUMxa9_and_b4), .B0(n3149), 
        .B1(output_p1_times_a1_mul_componentxUMxa11_and_b2), .Y(n3150) );
  NOR2X1 U2736 ( .A(n4528), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b10) );
  NOR2X1 U2737 ( .A(n4527), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b11) );
  NOR2X1 U2738 ( .A(n4527), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b11) );
  NOR2X1 U2739 ( .A(n4526), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b12) );
  NOR2X1 U2740 ( .A(n4526), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b12) );
  NOR2X1 U2741 ( .A(n231), .B(n4524), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b14) );
  NOR2X1 U2742 ( .A(n231), .B(n4523), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b15) );
  NOR2X1 U2743 ( .A(n213), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b8) );
  NOR2X1 U2744 ( .A(n214), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b7) );
  NOR2X1 U2745 ( .A(n213), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b8) );
  NOR2X1 U2746 ( .A(n212), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b9) );
  NOR2X1 U2747 ( .A(n214), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b7) );
  NOR2X1 U2748 ( .A(n213), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b8) );
  NOR2X1 U2749 ( .A(n212), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b9) );
  XOR2X1 U2750 ( .A(output_p1_times_a1_mul_componentxUMxa11_and_b2), .B(n3149), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127636032_127637936_127713632)
         );
  XOR2X1 U2751 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b6), .B(n3155), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732704_127722384_127724288)
         );
  XOR2X1 U2752 ( .A(output_p1_times_a1_mul_componentxUMxa12_and_b2), 
        .B(output_p1_times_a1_mul_componentxUMxa13_and_b1), .Y(n3159) );
  XOR2X1 U2753 ( .A(output_p1_times_a1_mul_componentxUMxa12_and_b3), 
        .B(output_p1_times_a1_mul_componentxUMxa13_and_b2), .Y(n3169) );
  XOR2X1 U2754 ( .A(output_p1_times_a1_mul_componentxUMxa15_and_b0), .B(n443), 
        .Y(n3231) );
  XOR2X1 U2755 ( .A(output_p1_times_a1_mul_componentxUMxa9_and_b4), 
        .B(output_p1_times_a1_mul_componentxUMxa10_and_b3), .Y(n3149) );
  XOR2X1 U2756 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b7), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b6), .Y(n3147) );
  XOR2X1 U2757 ( .A(output_p1_times_a1_mul_componentxUMxa9_and_b5), 
        .B(output_p1_times_a1_mul_componentxUMxa10_and_b4), .Y(n3157) );
  AND2X2 U2758 ( .A(output_p1_times_a1_mul_componentxUMxa13_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa12_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer1_127715536_127848576)
         );
  OR3XL U2759 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[1]), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[2]), 
        .C(output_p1_times_a1_mul_componentxUMxfirst_vector[0]), .Y(n3813) );
  XOR2X1 U2760 ( .A(output_p1_times_a1_mul_componentxUMxa14_and_b0), .B(n3159), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127715648_127848688_127850592)
         );
  XOR2X1 U2761 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b5), .B(n3147), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732592_127722272_127724176)
         );
  XOR2X1 U2762 ( .A(output_p1_times_a1_mul_componentxUMxa10_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa9_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127635696_127637600)
         );
  XOR2X1 U2763 ( .A(output_p1_times_a1_mul_componentxUMxa11_and_b1), .B(n3141), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127635920_127637824_127713520)
         );
  XOR2X1 U2764 ( .A(output_p1_times_a1_mul_componentxUMxa11_and_b3), .B(n3157), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127636144_127638048_127713744)
         );
  XOR2X1 U2765 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b1), .B(n3093), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127830448_127844704_127846608)
         );
  XOR2X1 U2766 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b6), .B(n3129), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127673344_127675248_127730464)
         );
  XOR2X1 U2767 ( .A(output_p1_times_a1_mul_componentxUMxa13_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa12_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127715536_127848576)
         );
  XOR2X1 U2768 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b3), .B(n3131), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127732368_127722048_127723952)
         );
  AND2X2 U2769 ( .A(output_p1_times_a1_mul_componentxUMxa10_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa9_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer1_127635696_127637600)
         );
  AND2X2 U2770 ( .A(output_p1_times_a1_mul_componentxUMxa1_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa0_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer1_127830168_127844480)
         );
  XOR2X1 U2771 ( .A(output_p1_times_a1_mul_componentxUMxa11_and_b0), .B(n3133), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127635808_127637712_127713408)
         );
  XOR2X1 U2772 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b0), .B(n3091), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127830336_127844592_127846496)
         );
  XOR2X1 U2773 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer4_128238312_128238424_128238592), 
        .B(n405), .Y(n3324) );
  XOR2X1 U2774 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer3_128264344_128264512), 
        .B(n3304), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer4_128238312_128238424_128238592)
         );
  INVX1 U2775 ( .A(n3318), .Y(n405) );
  XOR2X1 U2776 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer2_128199816_128200040_128199984), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer2_128199368_128199480_128199648), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer3_128264344_128264512)
         );
  INVX1 U2777 ( .A(n3158), .Y(n490) );
  AOI22X1 U2778 ( .A0(output_p1_times_a1_mul_componentxUMxa10_and_b4), 
        .A1(output_p1_times_a1_mul_componentxUMxa9_and_b5), .B0(n3157), 
        .B1(output_p1_times_a1_mul_componentxUMxa11_and_b3), .Y(n3158) );
  INVX1 U2779 ( .A(n3170), .Y(n507) );
  AOI22X1 U2780 ( .A0(output_p1_times_a1_mul_componentxUMxa13_and_b2), 
        .A1(output_p1_times_a1_mul_componentxUMxa12_and_b3), .B0(n3169), 
        .B1(output_p1_times_a1_mul_componentxUMxa14_and_b1), .Y(n3170) );
  INVX1 U2781 ( .A(n3156), .Y(n466) );
  AOI22X1 U2782 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b7), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b8), .B0(n3155), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b6), .Y(n3156) );
  INVX1 U2783 ( .A(n3160), .Y(n514) );
  AOI22X1 U2784 ( .A0(output_p1_times_a1_mul_componentxUMxa13_and_b1), 
        .A1(output_p1_times_a1_mul_componentxUMxa12_and_b2), .B0(n3159), 
        .B1(output_p1_times_a1_mul_componentxUMxa14_and_b0), .Y(n3160) );
  INVX1 U2785 ( .A(n3140), .Y(n485) );
  AOI22X1 U2786 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b5), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b6), .B0(n3139), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b4), .Y(n3140) );
  INVX1 U2787 ( .A(n3126), .Y(n499) );
  AOI22X1 U2788 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b3), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b4), .B0(n3125), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b2), .Y(n3126) );
  INVX1 U2789 ( .A(n3148), .Y(n474) );
  AOI22X1 U2790 ( .A0(output_p1_times_a1_mul_componentxUMxa7_and_b6), 
        .A1(output_p1_times_a1_mul_componentxUMxa6_and_b7), .B0(n3147), 
        .B1(output_p1_times_a1_mul_componentxUMxa8_and_b5), .Y(n3148) );
  NOR2X1 U2791 ( .A(n4526), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b12) );
  NOR2X1 U2792 ( .A(n4523), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b15) );
  NOR2X1 U2793 ( .A(n213), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b8) );
  NOR2X1 U2794 ( .A(n212), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b9) );
  NOR2X1 U2795 ( .A(n4528), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b10) );
  INVX1 U2796 ( .A(n3168), .Y(n484) );
  AOI22X1 U2797 ( .A0(output_p1_times_a1_mul_componentxUMxa10_and_b5), 
        .A1(output_p1_times_a1_mul_componentxUMxa9_and_b6), .B0(n3167), 
        .B1(output_p1_times_a1_mul_componentxUMxa11_and_b4), .Y(n3168) );
  AOI22X1 U2798 ( .A0(output_p1_times_a1_mul_componentxUMxa13_and_b3), 
        .A1(output_p1_times_a1_mul_componentxUMxa12_and_b4), .B0(n3179), 
        .B1(output_p1_times_a1_mul_componentxUMxa14_and_b2), .Y(n3180) );
  NOR2X1 U2799 ( .A(n4528), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b10) );
  NOR2X1 U2800 ( .A(n4527), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b11) );
  NOR2X1 U2801 ( .A(n4525), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b13) );
  NOR2X1 U2802 ( .A(n4525), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b13) );
  NOR2X1 U2803 ( .A(n4524), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b14) );
  NOR2X1 U2804 ( .A(n231), .B(n4522), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b16) );
  XOR2X1 U2805 ( .A(output_p1_times_a1_mul_componentxUMxa1_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa0_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[1]) );
  NOR2X1 U2806 ( .A(n212), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b9) );
  NOR2X1 U2807 ( .A(n222), .B(n214), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b7) );
  NOR2X1 U2808 ( .A(n214), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b7) );
  NOR2X1 U2809 ( .A(n213), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b8) );
  NOR2X1 U2810 ( .A(n214), .B(n4545), 
        .Y(output_p1_times_a1_mul_componentxUMxa10_and_b7) );
  NOR2X1 U2811 ( .A(n4525), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b13) );
  NOR2X1 U2812 ( .A(n4522), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b16) );
  XOR2X1 U2813 ( .A(output_p1_times_a1_mul_componentxUMxa12_and_b4), 
        .B(output_p1_times_a1_mul_componentxUMxa13_and_b3), .Y(n3179) );
  XOR2X1 U2814 ( .A(output_p1_times_a1_mul_componentxUMxa9_and_b6), 
        .B(output_p1_times_a1_mul_componentxUMxa10_and_b5), .Y(n3167) );
  XOR2X1 U2815 ( .A(output_p1_times_a1_mul_componentxUMxa9_and_b7), 
        .B(output_p1_times_a1_mul_componentxUMxa10_and_b6), .Y(n3177) );
  XOR2X1 U2816 ( .A(output_p1_times_a1_mul_componentxUMxa11_and_b5), .B(n3177), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127636368_127638272_127713968)
         );
  XOR2X1 U2817 ( .A(output_p1_times_a1_mul_componentxUMxa11_and_b4), .B(n3167), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127636256_127638160_127713856)
         );
  XOR2X1 U2818 ( .A(output_p1_times_a1_mul_componentxUMxa14_and_b2), .B(n3179), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127715872_127848912_127850816)
         );
  XOR2X1 U2819 ( .A(output_p1_times_a1_mul_componentxUMxa14_and_b1), .B(n3169), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127715760_127848800_127850704)
         );
  XOR2X1 U2820 ( .A(output_p1_times_a1_mul_componentxUMxa16_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa15_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127627504_127629408)
         );
  XOR2X1 U2821 ( .A(output_p1_times_a1_mul_componentxUMxa5_and_b12), .B(n3182), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127674016_127675920_127731136)
         );
  NOR2X1 U2822 ( .A(n4526), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b12) );
  XOR2X1 U2823 ( .A(output_p1_times_a1_mul_componentxUMxa3_and_b14), 
        .B(output_p1_times_a1_mul_componentxUMxa4_and_b13), .Y(n3182) );
  NOR2X1 U2824 ( .A(n4524), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b14) );
  XOR2X1 U2825 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127733040_127722720_127724624), 
        .B(n3245), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128199368_128199480_128199648)
         );
  XOR2X1 U2826 ( .A(output_p1_times_a1_mul_componentxUMxa8_and_b9), .B(n3183), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127733040_127722720_127724624)
         );
  XOR2X1 U2827 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127832016_127846272_127848176), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127674016_127675920_127731136), 
        .Y(n3245) );
  NOR2X1 U2828 ( .A(n212), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b9) );
  XOR2X1 U2829 ( .A(n3178), .B(n3180), .Y(n3244) );
  AOI22X1 U2830 ( .A0(output_p1_times_a1_mul_componentxUMxa10_and_b6), 
        .A1(output_p1_times_a1_mul_componentxUMxa9_and_b7), .B0(n3177), 
        .B1(output_p1_times_a1_mul_componentxUMxa11_and_b5), .Y(n3178) );
  INVX1 U2831 ( .A(n4555), .Y(n516) );
  AOI22XL U2832 ( .A0(output_p1_times_a1_mul_componentxUMxfirst_vector[2]), 
        .A1(n113), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[2]), 
        .B1(n4548), .Y(n4555) );
  XNOR2X1 U2833 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[2]), 
        .B(n3814), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[2]) );
  NOR2X1 U2834 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[0]), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[1]), .Y(n3814) );
  INVX1 U2835 ( .A(n4556), .Y(n517) );
  AOI22XL U2836 ( .A0(output_p1_times_a1_mul_componentxUMxfirst_vector[1]), 
        .A1(n114), 
        .B0(output_p1_times_a1_mul_componentxunsigned_output_inverted[1]), 
        .B1(n4548), .Y(n4556) );
  XOR2X1 U2837 ( .A(output_p1_times_a1_mul_componentxUMxfirst_vector[1]), 
        .B(output_p1_times_a1_mul_componentxUMxfirst_vector[0]), 
        .Y(output_p1_times_a1_mul_componentxunsigned_output_inverted[1]) );
  XOR2X1 U2838 ( .A(output_p1_times_a1_mul_componentxUMxa2_and_b15), .B(n3181), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127832016_127846272_127848176)
         );
  NOR2X1 U2839 ( .A(n4523), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b15) );
  XOR2X1 U2840 ( .A(output_p1_times_a1_mul_componentxUMxa0_and_b17), 
        .B(output_p1_times_a1_mul_componentxUMxa1_and_b16), .Y(n3181) );
  NOR2X1 U2841 ( .A(n231), .B(n20), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b17) );
  INVX1 U2842 ( .A(n3232), .Y(n410) );
  AOI22X1 U2843 ( .A0(n443), 
        .A1(output_p1_times_a1_mul_componentxUMxa15_and_b0), .B0(n3231), 
        .B1(n411), .Y(n3232) );
  AND2X2 U2844 ( .A(output_p1_times_a1_mul_componentxUMxa16_and_b0), 
        .B(output_p1_times_a1_mul_componentxUMxa15_and_b1), 
        .Y(output_p1_times_a1_mul_componentxUMxcarry_layer1_127627504_127629408)
         );
  INVX1 U2845 ( .A(n4565), .Y(n518) );
  AOI22XL U2846 ( .A0(output_p1_times_a1_mul_componentxUMxfirst_vector[0]), 
        .A1(n113), .B0(output_p1_times_a1_mul_componentxUMxfirst_vector[0]), 
        .B1(n4548), .Y(n4565) );
  XOR2X1 U2847 ( .A(output_p1_times_a1_mul_componentxUMxa6_and_b11), 
        .B(output_p1_times_a1_mul_componentxUMxa7_and_b10), .Y(n3183) );
  NOR2X1 U2848 ( .A(n4527), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b11) );
  NOR2X1 U2849 ( .A(n4528), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b10) );
  XOR2X1 U2850 ( .A(n134), .B(n361), .Y(n80) );
  INVX1 U2851 ( .A(n80), .Y(n4548) );
  XOR2X1 U2852 ( .A(input_p1_times_b1_mul_componentxUMxa9_and_b2), 
        .B(input_p1_times_b1_mul_componentxUMxa10_and_b1), .Y(n2665) );
  XOR2X1 U2853 ( .A(input_p2_times_b2_mul_componentxUMxa9_and_b2), 
        .B(input_p2_times_b2_mul_componentxUMxa10_and_b1), .Y(n2899) );
  XOR2X1 U2854 ( .A(output_p2_times_a2_mul_componentxUMxa9_and_b2), 
        .B(output_p2_times_a2_mul_componentxUMxa10_and_b1), .Y(n3367) );
  XOR2X1 U2855 ( .A(input_times_b0_mul_componentxUMxa9_and_b2), 
        .B(input_times_b0_mul_componentxUMxa10_and_b1), .Y(n2431) );
  INVX1 U2856 ( .A(n2666), .Y(n988) );
  AOI22X1 U2857 ( .A0(input_p1_times_b1_mul_componentxUMxa10_and_b1), 
        .A1(input_p1_times_b1_mul_componentxUMxa9_and_b2), .B0(n2665), 
        .B1(input_p1_times_b1_mul_componentxUMxa11_and_b0), .Y(n2666) );
  INVX1 U2858 ( .A(n2900), .Y(n1147) );
  AOI22X1 U2859 ( .A0(input_p2_times_b2_mul_componentxUMxa10_and_b1), 
        .A1(input_p2_times_b2_mul_componentxUMxa9_and_b2), .B0(n2899), 
        .B1(input_p2_times_b2_mul_componentxUMxa11_and_b0), .Y(n2900) );
  INVX1 U2860 ( .A(n3368), .Y(n670) );
  AOI22X1 U2861 ( .A0(output_p2_times_a2_mul_componentxUMxa10_and_b1), 
        .A1(output_p2_times_a2_mul_componentxUMxa9_and_b2), .B0(n3367), 
        .B1(output_p2_times_a2_mul_componentxUMxa11_and_b0), .Y(n3368) );
  INVX1 U2862 ( .A(n2432), .Y(n829) );
  AOI22X1 U2863 ( .A0(input_times_b0_mul_componentxUMxa10_and_b1), 
        .A1(input_times_b0_mul_componentxUMxa9_and_b2), .B0(n2431), 
        .B1(input_times_b0_mul_componentxUMxa11_and_b0), .Y(n2432) );
  INVX1 U2864 ( .A(n2674), .Y(n981) );
  AOI22X1 U2865 ( .A0(input_p1_times_b1_mul_componentxUMxa10_and_b2), 
        .A1(input_p1_times_b1_mul_componentxUMxa9_and_b3), .B0(n2673), 
        .B1(input_p1_times_b1_mul_componentxUMxa11_and_b1), .Y(n2674) );
  INVX1 U2866 ( .A(n2440), .Y(n822) );
  AOI22X1 U2867 ( .A0(input_times_b0_mul_componentxUMxa10_and_b2), 
        .A1(input_times_b0_mul_componentxUMxa9_and_b3), .B0(n2439), 
        .B1(input_times_b0_mul_componentxUMxa11_and_b1), .Y(n2440) );
  INVX1 U2868 ( .A(n2682), .Y(n975) );
  AOI22X1 U2869 ( .A0(input_p1_times_b1_mul_componentxUMxa10_and_b3), 
        .A1(input_p1_times_b1_mul_componentxUMxa9_and_b4), .B0(n2681), 
        .B1(input_p1_times_b1_mul_componentxUMxa11_and_b2), .Y(n2682) );
  INVX1 U2870 ( .A(n2448), .Y(n816) );
  AOI22X1 U2871 ( .A0(input_times_b0_mul_componentxUMxa10_and_b3), 
        .A1(input_times_b0_mul_componentxUMxa9_and_b4), .B0(n2447), 
        .B1(input_times_b0_mul_componentxUMxa11_and_b2), .Y(n2448) );
  INVX1 U2872 ( .A(n2628), .Y(n978) );
  AOI22X1 U2873 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b3), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b4), .B0(n2627), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b2), .Y(n2628) );
  INVX1 U2874 ( .A(n2862), .Y(n1137) );
  AOI22X1 U2875 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b3), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b4), .B0(n2861), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b2), .Y(n2862) );
  INVX1 U2876 ( .A(n3330), .Y(n660) );
  AOI22X1 U2877 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b3), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b4), .B0(n3329), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b2), .Y(n3330) );
  INVX1 U2878 ( .A(n2394), .Y(n819) );
  AOI22X1 U2879 ( .A0(input_times_b0_mul_componentxUMxa1_and_b3), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b4), .B0(n2393), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b2), .Y(n2394) );
  INVX1 U2880 ( .A(n2630), .Y(n971) );
  AOI22X1 U2881 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b4), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b5), .B0(n2629), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b3), .Y(n2630) );
  INVX1 U2882 ( .A(n2396), .Y(n812) );
  AOI22X1 U2883 ( .A0(input_times_b0_mul_componentxUMxa1_and_b4), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b5), .B0(n2395), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b3), .Y(n2396) );
  INVX1 U2884 ( .A(n2860), .Y(n1144) );
  AOI22X1 U2885 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b2), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b3), .B0(n2859), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b1), .Y(n2860) );
  INVX1 U2886 ( .A(n3328), .Y(n667) );
  AOI22X1 U2887 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b2), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b3), .B0(n3327), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b1), .Y(n3328) );
  INVX1 U2888 ( .A(n2636), .Y(n983) );
  AOI22X1 U2889 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b2), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b3), .B0(n2635), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b1), .Y(n2636) );
  INVX1 U2890 ( .A(n2874), .Y(n1136) );
  AOI22X1 U2891 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b3), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b4), .B0(n2873), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b2), .Y(n2874) );
  INVX1 U2892 ( .A(n2872), .Y(n1115) );
  AOI22X1 U2893 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b6), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b7), .B0(n2871), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b5), .Y(n2872) );
  INVX1 U2894 ( .A(n3342), .Y(n659) );
  AOI22X1 U2895 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b3), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b4), .B0(n3341), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b2), .Y(n3342) );
  INVX1 U2896 ( .A(n3340), .Y(n638) );
  AOI22X1 U2897 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b6), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b7), .B0(n3339), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b5), .Y(n3340) );
  INVX1 U2898 ( .A(n2402), .Y(n824) );
  AOI22X1 U2899 ( .A0(input_times_b0_mul_componentxUMxa4_and_b2), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b3), .B0(n2401), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b1), .Y(n2402) );
  INVX1 U2900 ( .A(n2726), .Y(n970) );
  AOI22X1 U2901 ( .A0(n971), .A1(input_p1_times_b1_mul_componentxUMxa6_and_b0), 
        .B0(n2725), .B1(n990), .Y(n2726) );
  INVX1 U2902 ( .A(n2646), .Y(n989) );
  AOI22X1 U2903 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b1), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b2), .B0(n2645), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b0), .Y(n2646) );
  INVX1 U2904 ( .A(n2960), .Y(n1129) );
  AOI22X1 U2905 ( .A0(n1130), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b0), .B0(n2959), 
        .B1(n1149), .Y(n2960) );
  INVX1 U2906 ( .A(n3428), .Y(n652) );
  AOI22X1 U2907 ( .A0(n653), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b0), .B0(n3427), 
        .B1(n672), .Y(n3428) );
  INVX1 U2908 ( .A(n2492), .Y(n811) );
  AOI22X1 U2909 ( .A0(n812), .A1(input_times_b0_mul_componentxUMxa6_and_b0), 
        .B0(n2491), .B1(n831), .Y(n2492) );
  INVX1 U2910 ( .A(n2412), .Y(n830) );
  AOI22X1 U2911 ( .A0(input_times_b0_mul_componentxUMxa7_and_b1), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b2), .B0(n2411), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b0), .Y(n2412) );
  INVX1 U2912 ( .A(n2734), .Y(n945) );
  AOI22X1 U2913 ( .A0(n946), .A1(input_p1_times_b1_mul_componentxUMxa9_and_b0), 
        .B0(n2733), .B1(n969), .Y(n2734) );
  INVX1 U2914 ( .A(n2664), .Y(n968) );
  AOI22X1 U2915 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b4), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b5), .B0(n2663), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b3), .Y(n2664) );
  INVX1 U2916 ( .A(n2898), .Y(n1127) );
  AOI22X1 U2917 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b4), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b5), .B0(n2897), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b3), .Y(n2898) );
  INVX1 U2918 ( .A(n3366), .Y(n650) );
  AOI22X1 U2919 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b4), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b5), .B0(n3365), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b3), .Y(n3366) );
  INVX1 U2920 ( .A(n2500), .Y(n786) );
  AOI22X1 U2921 ( .A0(n787), .A1(input_times_b0_mul_componentxUMxa9_and_b0), 
        .B0(n2499), .B1(n810), .Y(n2500) );
  INVX1 U2922 ( .A(n2430), .Y(n809) );
  AOI22X1 U2923 ( .A0(input_times_b0_mul_componentxUMxa7_and_b4), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b5), .B0(n2429), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b3), .Y(n2430) );
  INVX1 U2924 ( .A(n2656), .Y(n953) );
  AOI22X1 U2925 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b6), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b7), .B0(n2655), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b5), .Y(n2656) );
  INVX1 U2926 ( .A(n2422), .Y(n794) );
  AOI22X1 U2927 ( .A0(input_times_b0_mul_componentxUMxa4_and_b6), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b7), .B0(n2421), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b5), .Y(n2422) );
  XOR2X1 U2928 ( .A(input_p1_times_b1_mul_componentxUMxa11_and_b2), .B(n2681), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127636032_127637936_127713632)
         );
  XOR2X1 U2929 ( .A(input_times_b0_mul_componentxUMxa11_and_b2), .B(n2447), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127636032_127637936_127713632)
         );
  XOR2X1 U2930 ( .A(input_p2_times_b2_mul_componentxUMxa11_and_b2), .B(n2915), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127636032_127637936_127713632)
         );
  XOR2X1 U2931 ( .A(output_p2_times_a2_mul_componentxUMxa11_and_b2), .B(n3383), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127636032_127637936_127713632)
         );
  XOR2X1 U2932 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b2), .B(n2627), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127830560_127844816_127846720)
         );
  XOR2X1 U2933 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b2), .B(n2861), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127830560_127844816_127846720)
         );
  XOR2X1 U2934 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b2), .B(n3329), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127830560_127844816_127846720)
         );
  XOR2X1 U2935 ( .A(input_times_b0_mul_componentxUMxa2_and_b2), .B(n2393), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127830560_127844816_127846720)
         );
  XOR2X1 U2936 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b3), .B(n2643), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673008_127674912_127730128)
         );
  XOR2X1 U2937 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b3), .B(n2877), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673008_127674912_127730128)
         );
  XOR2X1 U2938 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b3), .B(n3345), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673008_127674912_127730128)
         );
  XOR2X1 U2939 ( .A(input_times_b0_mul_componentxUMxa5_and_b3), .B(n2409), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673008_127674912_127730128)
         );
  XOR2X1 U2940 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b4), .B(n2671), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732480_127722160_127724064)
         );
  XOR2X1 U2941 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b4), .B(n2905), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732480_127722160_127724064)
         );
  XOR2X1 U2942 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b4), .B(n3373), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732480_127722160_127724064)
         );
  XOR2X1 U2943 ( .A(input_times_b0_mul_componentxUMxa8_and_b4), .B(n2437), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732480_127722160_127724064)
         );
  XOR2X1 U2944 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b5), .B(n2655), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673232_127675136_127730352)
         );
  XOR2X1 U2945 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b5), .B(n2889), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673232_127675136_127730352)
         );
  XOR2X1 U2946 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b5), .B(n3357), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673232_127675136_127730352)
         );
  XOR2X1 U2947 ( .A(input_times_b0_mul_componentxUMxa5_and_b5), .B(n2421), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673232_127675136_127730352)
         );
  XOR2X1 U2948 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b6), .B(n2687), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732704_127722384_127724288)
         );
  XOR2X1 U2949 ( .A(input_times_b0_mul_componentxUMxa8_and_b6), .B(n2453), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732704_127722384_127724288)
         );
  XOR2X1 U2950 ( .A(input_p1_times_b1_mul_componentxUMxa12_and_b0), .B(n912), 
        .Y(n2745) );
  XOR2X1 U2951 ( .A(input_times_b0_mul_componentxUMxa12_and_b0), .B(n753), 
        .Y(n2511) );
  XOR2X1 U2952 ( .A(input_p1_times_b1_mul_componentxUMxa12_and_b2), 
        .B(input_p1_times_b1_mul_componentxUMxa13_and_b1), .Y(n2691) );
  XOR2X1 U2953 ( .A(input_times_b0_mul_componentxUMxa12_and_b2), 
        .B(input_times_b0_mul_componentxUMxa13_and_b1), .Y(n2457) );
  XOR2X1 U2954 ( .A(input_p1_times_b1_mul_componentxUMxa12_and_b3), 
        .B(input_p1_times_b1_mul_componentxUMxa13_and_b2), .Y(n2701) );
  XOR2X1 U2955 ( .A(input_times_b0_mul_componentxUMxa12_and_b3), 
        .B(input_times_b0_mul_componentxUMxa13_and_b2), .Y(n2467) );
  XOR2X1 U2956 ( .A(input_p2_times_b2_mul_componentxUMxa12_and_b0), .B(n1071), 
        .Y(n2979) );
  XOR2X1 U2957 ( .A(output_p2_times_a2_mul_componentxUMxa12_and_b0), .B(n594), 
        .Y(n3447) );
  XOR2X1 U2958 ( .A(input_p2_times_b2_mul_componentxUMxa12_and_b2), 
        .B(input_p2_times_b2_mul_componentxUMxa13_and_b1), .Y(n2925) );
  XOR2X1 U2959 ( .A(output_p2_times_a2_mul_componentxUMxa12_and_b2), 
        .B(output_p2_times_a2_mul_componentxUMxa13_and_b1), .Y(n3393) );
  XOR2X1 U2960 ( .A(input_p2_times_b2_mul_componentxUMxa12_and_b3), 
        .B(input_p2_times_b2_mul_componentxUMxa13_and_b2), .Y(n2935) );
  XOR2X1 U2961 ( .A(output_p2_times_a2_mul_componentxUMxa12_and_b3), 
        .B(output_p2_times_a2_mul_componentxUMxa13_and_b2), .Y(n3403) );
  XOR2X1 U2962 ( .A(input_p1_times_b1_mul_componentxUMxa15_and_b0), .B(n919), 
        .Y(n2763) );
  XOR2X1 U2963 ( .A(input_times_b0_mul_componentxUMxa15_and_b0), .B(n760), 
        .Y(n2529) );
  XOR2X1 U2964 ( .A(input_p2_times_b2_mul_componentxUMxa15_and_b0), .B(n1078), 
        .Y(n2997) );
  XOR2X1 U2965 ( .A(output_p2_times_a2_mul_componentxUMxa15_and_b0), .B(n601), 
        .Y(n3465) );
  XOR2X1 U2966 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b4), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b3), .Y(n2627) );
  XOR2X1 U2967 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b4), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b3), .Y(n2861) );
  XOR2X1 U2968 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b4), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b3), .Y(n3329) );
  XOR2X1 U2969 ( .A(input_times_b0_mul_componentxUMxa0_and_b4), 
        .B(input_times_b0_mul_componentxUMxa1_and_b3), .Y(n2393) );
  XOR2X1 U2970 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b5), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b4), .Y(n2629) );
  XOR2X1 U2971 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b5), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b4), .Y(n2863) );
  XOR2X1 U2972 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b5), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b4), .Y(n3331) );
  XOR2X1 U2973 ( .A(input_times_b0_mul_componentxUMxa0_and_b5), 
        .B(input_times_b0_mul_componentxUMxa1_and_b4), .Y(n2395) );
  XOR2X1 U2974 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b3), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b2), .Y(n2625) );
  XOR2X1 U2975 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b3), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b2), .Y(n2859) );
  XOR2X1 U2976 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b3), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b2), .Y(n3327) );
  XOR2X1 U2977 ( .A(input_times_b0_mul_componentxUMxa0_and_b3), 
        .B(input_times_b0_mul_componentxUMxa1_and_b2), .Y(n2391) );
  XOR2X1 U2978 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b8), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b7), .Y(n2641) );
  XOR2X1 U2979 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b7), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b6), .Y(n2637) );
  XOR2X1 U2980 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b8), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b7), .Y(n2875) );
  XOR2X1 U2981 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b7), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b6), .Y(n2871) );
  XOR2X1 U2982 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b8), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b7), .Y(n3343) );
  XOR2X1 U2983 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b7), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b6), .Y(n3339) );
  XOR2X1 U2984 ( .A(input_times_b0_mul_componentxUMxa0_and_b8), 
        .B(input_times_b0_mul_componentxUMxa1_and_b7), .Y(n2407) );
  XOR2X1 U2985 ( .A(input_times_b0_mul_componentxUMxa0_and_b7), 
        .B(input_times_b0_mul_componentxUMxa1_and_b6), .Y(n2403) );
  XOR2X1 U2986 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b0), .B(n971), 
        .Y(n2725) );
  XOR2X1 U2987 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b6), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b5), .Y(n2633) );
  XOR2X1 U2988 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b0), .B(n1130), 
        .Y(n2959) );
  XOR2X1 U2989 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b6), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b5), .Y(n2867) );
  XOR2X1 U2990 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b0), .B(n653), 
        .Y(n3427) );
  XOR2X1 U2991 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b6), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b5), .Y(n3335) );
  XOR2X1 U2992 ( .A(input_times_b0_mul_componentxUMxa6_and_b0), .B(n812), 
        .Y(n2491) );
  XOR2X1 U2993 ( .A(input_times_b0_mul_componentxUMxa0_and_b6), 
        .B(input_times_b0_mul_componentxUMxa1_and_b5), .Y(n2399) );
  XOR2X1 U2994 ( .A(input_p1_times_b1_mul_componentxUMxa9_and_b0), .B(n946), 
        .Y(n2733) );
  XOR2X1 U2995 ( .A(input_p2_times_b2_mul_componentxUMxa9_and_b0), .B(n1105), 
        .Y(n2967) );
  XOR2X1 U2996 ( .A(output_p2_times_a2_mul_componentxUMxa9_and_b0), .B(n628), 
        .Y(n3435) );
  XOR2X1 U2997 ( .A(input_times_b0_mul_componentxUMxa9_and_b0), .B(n787), 
        .Y(n2499) );
  XOR2X1 U2998 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b2), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b1), .Y(n2631) );
  XOR2X1 U2999 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b2), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b1), .Y(n2865) );
  XOR2X1 U3000 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b2), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b1), .Y(n3333) );
  XOR2X1 U3001 ( .A(input_times_b0_mul_componentxUMxa3_and_b2), 
        .B(input_times_b0_mul_componentxUMxa4_and_b1), .Y(n2397) );
  XOR2X1 U3002 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b2), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b1), .Y(n2645) );
  XOR2X1 U3003 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b2), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b1), .Y(n2879) );
  XOR2X1 U3004 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b2), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b1), .Y(n3347) );
  XOR2X1 U3005 ( .A(input_times_b0_mul_componentxUMxa6_and_b2), 
        .B(input_times_b0_mul_componentxUMxa7_and_b1), .Y(n2411) );
  XOR2X1 U3006 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b3), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b2), .Y(n2635) );
  XOR2X1 U3007 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b3), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b2), .Y(n2869) );
  XOR2X1 U3008 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b3), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b2), .Y(n3337) );
  XOR2X1 U3009 ( .A(input_times_b0_mul_componentxUMxa3_and_b3), 
        .B(input_times_b0_mul_componentxUMxa4_and_b2), .Y(n2401) );
  XOR2X1 U3010 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b3), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b2), .Y(n2651) );
  XOR2X1 U3011 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b3), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b2), .Y(n2885) );
  XOR2X1 U3012 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b3), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b2), .Y(n3353) );
  XOR2X1 U3013 ( .A(input_times_b0_mul_componentxUMxa6_and_b3), 
        .B(input_times_b0_mul_componentxUMxa7_and_b2), .Y(n2417) );
  XOR2X1 U3014 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b4), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b3), .Y(n2639) );
  XOR2X1 U3015 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b4), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b3), .Y(n2873) );
  XOR2X1 U3016 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b4), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b3), .Y(n3341) );
  XOR2X1 U3017 ( .A(input_times_b0_mul_componentxUMxa3_and_b4), 
        .B(input_times_b0_mul_componentxUMxa4_and_b3), .Y(n2405) );
  XOR2X1 U3018 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b4), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b3), .Y(n2657) );
  XOR2X1 U3019 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b4), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b3), .Y(n2891) );
  XOR2X1 U3020 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b4), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b3), .Y(n3359) );
  XOR2X1 U3021 ( .A(input_times_b0_mul_componentxUMxa6_and_b4), 
        .B(input_times_b0_mul_componentxUMxa7_and_b3), .Y(n2423) );
  XOR2X1 U3022 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b5), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b4), .Y(n2643) );
  XOR2X1 U3023 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b5), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b4), .Y(n2877) );
  XOR2X1 U3024 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b5), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b4), .Y(n3345) );
  XOR2X1 U3025 ( .A(input_times_b0_mul_componentxUMxa3_and_b5), 
        .B(input_times_b0_mul_componentxUMxa4_and_b4), .Y(n2409) );
  XOR2X1 U3026 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b5), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b4), .Y(n2663) );
  XOR2X1 U3027 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b5), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b4), .Y(n2897) );
  XOR2X1 U3028 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b5), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b4), .Y(n3365) );
  XOR2X1 U3029 ( .A(input_times_b0_mul_componentxUMxa6_and_b5), 
        .B(input_times_b0_mul_componentxUMxa7_and_b4), .Y(n2429) );
  XOR2X1 U3030 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b6), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b5), .Y(n2649) );
  XOR2X1 U3031 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b6), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b5), .Y(n2883) );
  XOR2X1 U3032 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b6), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b5), .Y(n3351) );
  XOR2X1 U3033 ( .A(input_times_b0_mul_componentxUMxa3_and_b6), 
        .B(input_times_b0_mul_componentxUMxa4_and_b5), .Y(n2415) );
  XOR2X1 U3034 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b6), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b5), .Y(n2671) );
  XOR2X1 U3035 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b6), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b5), .Y(n2905) );
  XOR2X1 U3036 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b6), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b5), .Y(n3373) );
  XOR2X1 U3037 ( .A(input_times_b0_mul_componentxUMxa6_and_b6), 
        .B(input_times_b0_mul_componentxUMxa7_and_b5), .Y(n2437) );
  XOR2X1 U3038 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b7), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b6), .Y(n2655) );
  XOR2X1 U3039 ( .A(input_p1_times_b1_mul_componentxUMxa9_and_b3), 
        .B(input_p1_times_b1_mul_componentxUMxa10_and_b2), .Y(n2673) );
  XOR2X1 U3040 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b7), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b6), .Y(n2889) );
  XOR2X1 U3041 ( .A(input_p2_times_b2_mul_componentxUMxa9_and_b3), 
        .B(input_p2_times_b2_mul_componentxUMxa10_and_b2), .Y(n2907) );
  XOR2X1 U3042 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b7), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b6), .Y(n3357) );
  XOR2X1 U3043 ( .A(output_p2_times_a2_mul_componentxUMxa9_and_b3), 
        .B(output_p2_times_a2_mul_componentxUMxa10_and_b2), .Y(n3375) );
  XOR2X1 U3044 ( .A(input_times_b0_mul_componentxUMxa3_and_b7), 
        .B(input_times_b0_mul_componentxUMxa4_and_b6), .Y(n2421) );
  XOR2X1 U3045 ( .A(input_times_b0_mul_componentxUMxa9_and_b3), 
        .B(input_times_b0_mul_componentxUMxa10_and_b2), .Y(n2439) );
  XOR2X1 U3046 ( .A(input_p1_times_b1_mul_componentxUMxa9_and_b4), 
        .B(input_p1_times_b1_mul_componentxUMxa10_and_b3), .Y(n2681) );
  XOR2X1 U3047 ( .A(input_p2_times_b2_mul_componentxUMxa9_and_b4), 
        .B(input_p2_times_b2_mul_componentxUMxa10_and_b3), .Y(n2915) );
  XOR2X1 U3048 ( .A(output_p2_times_a2_mul_componentxUMxa9_and_b4), 
        .B(output_p2_times_a2_mul_componentxUMxa10_and_b3), .Y(n3383) );
  XOR2X1 U3049 ( .A(input_times_b0_mul_componentxUMxa9_and_b4), 
        .B(input_times_b0_mul_componentxUMxa10_and_b3), .Y(n2447) );
  XOR2X1 U3050 ( .A(input_p1_times_b1_mul_componentxUMxa9_and_b5), 
        .B(input_p1_times_b1_mul_componentxUMxa10_and_b4), .Y(n2689) );
  XOR2X1 U3051 ( .A(input_p2_times_b2_mul_componentxUMxa9_and_b5), 
        .B(input_p2_times_b2_mul_componentxUMxa10_and_b4), .Y(n2923) );
  XOR2X1 U3052 ( .A(output_p2_times_a2_mul_componentxUMxa9_and_b5), 
        .B(output_p2_times_a2_mul_componentxUMxa10_and_b4), .Y(n3391) );
  XOR2X1 U3053 ( .A(input_times_b0_mul_componentxUMxa9_and_b5), 
        .B(input_times_b0_mul_componentxUMxa10_and_b4), .Y(n2455) );
  XOR2X1 U3054 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b8), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b7), .Y(n2687) );
  XOR2X1 U3055 ( .A(input_times_b0_mul_componentxUMxa6_and_b8), 
        .B(input_times_b0_mul_componentxUMxa7_and_b7), .Y(n2453) );
  AND2X2 U3056 ( .A(input_p1_times_b1_mul_componentxUMxa13_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa12_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer1_127715536_127848576)
         );
  AND2X2 U3057 ( .A(input_times_b0_mul_componentxUMxa13_and_b0), 
        .B(input_times_b0_mul_componentxUMxa12_and_b1), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer1_127715536_127848576)
         );
  AND2X2 U3058 ( .A(input_p2_times_b2_mul_componentxUMxa13_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa12_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer1_127715536_127848576)
         );
  AND2X2 U3059 ( .A(output_p2_times_a2_mul_componentxUMxa13_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa12_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer1_127715536_127848576)
         );
  AND2X2 U3060 ( .A(input_p1_times_b1_mul_componentxUMxa4_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa3_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer1_127672560_127674464)
         );
  AND2X2 U3061 ( .A(input_p2_times_b2_mul_componentxUMxa4_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa3_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer1_127672560_127674464)
         );
  AND2X2 U3062 ( .A(output_p2_times_a2_mul_componentxUMxa4_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa3_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer1_127672560_127674464)
         );
  AND2X2 U3063 ( .A(input_times_b0_mul_componentxUMxa4_and_b0), 
        .B(input_times_b0_mul_componentxUMxa3_and_b1), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer1_127672560_127674464)
         );
  XOR2X1 U3064 ( .A(input_p1_times_b1_mul_componentxUMxa14_and_b0), .B(n2691), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127715648_127848688_127850592)
         );
  XOR2X1 U3065 ( .A(input_times_b0_mul_componentxUMxa14_and_b0), .B(n2457), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127715648_127848688_127850592)
         );
  XOR2X1 U3066 ( .A(input_p2_times_b2_mul_componentxUMxa14_and_b0), .B(n2925), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127715648_127848688_127850592)
         );
  XOR2X1 U3067 ( .A(output_p2_times_a2_mul_componentxUMxa14_and_b0), .B(n3393), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127715648_127848688_127850592)
         );
  XOR2X1 U3068 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b1), .B(n2651), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732144_127721824_127723728)
         );
  XOR2X1 U3069 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b1), .B(n2885), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732144_127721824_127723728)
         );
  XOR2X1 U3070 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b1), .B(n3353), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732144_127721824_127723728)
         );
  XOR2X1 U3071 ( .A(input_times_b0_mul_componentxUMxa8_and_b1), .B(n2417), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732144_127721824_127723728)
         );
  XOR2X1 U3072 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b6), .B(n2641), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831008_127845264_127847168)
         );
  XOR2X1 U3073 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b6), .B(n2875), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831008_127845264_127847168)
         );
  XOR2X1 U3074 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b6), .B(n3343), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831008_127845264_127847168)
         );
  XOR2X1 U3075 ( .A(input_times_b0_mul_componentxUMxa2_and_b6), .B(n2407), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831008_127845264_127847168)
         );
  XOR2X1 U3076 ( .A(input_p1_times_b1_mul_componentxUMxa10_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa9_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127635696_127637600)
         );
  XOR2X1 U3077 ( .A(input_p2_times_b2_mul_componentxUMxa10_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa9_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127635696_127637600)
         );
  XOR2X1 U3078 ( .A(output_p2_times_a2_mul_componentxUMxa10_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa9_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127635696_127637600)
         );
  XOR2X1 U3079 ( .A(input_times_b0_mul_componentxUMxa10_and_b0), 
        .B(input_times_b0_mul_componentxUMxa9_and_b1), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127635696_127637600) );
  XOR2X1 U3080 ( .A(input_p1_times_b1_mul_componentxUMxa11_and_b1), .B(n2673), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127635920_127637824_127713520)
         );
  XOR2X1 U3081 ( .A(input_times_b0_mul_componentxUMxa11_and_b1), .B(n2439), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127635920_127637824_127713520)
         );
  XOR2X1 U3082 ( .A(input_p1_times_b1_mul_componentxUMxa11_and_b3), .B(n2689), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127636144_127638048_127713744)
         );
  XOR2X1 U3083 ( .A(input_times_b0_mul_componentxUMxa11_and_b3), .B(n2455), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127636144_127638048_127713744)
         );
  XOR2X1 U3084 ( .A(input_p2_times_b2_mul_componentxUMxa11_and_b1), .B(n2907), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127635920_127637824_127713520)
         );
  XOR2X1 U3085 ( .A(output_p2_times_a2_mul_componentxUMxa11_and_b1), .B(n3375), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127635920_127637824_127713520)
         );
  XOR2X1 U3086 ( .A(input_p2_times_b2_mul_componentxUMxa11_and_b3), .B(n2923), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127636144_127638048_127713744)
         );
  XOR2X1 U3087 ( .A(output_p2_times_a2_mul_componentxUMxa11_and_b3), .B(n3391), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127636144_127638048_127713744)
         );
  XOR2X1 U3088 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b0), .B(n2645), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732032_127721712_127723616)
         );
  XOR2X1 U3089 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b0), .B(n2879), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732032_127721712_127723616)
         );
  XOR2X1 U3090 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b0), .B(n3347), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732032_127721712_127723616)
         );
  XOR2X1 U3091 ( .A(input_times_b0_mul_componentxUMxa8_and_b0), .B(n2411), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732032_127721712_127723616)
         );
  XOR2X1 U3092 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b2), .B(n2657), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732256_127721936_127723840)
         );
  XOR2X1 U3093 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b2), .B(n2891), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732256_127721936_127723840)
         );
  XOR2X1 U3094 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b2), .B(n3359), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732256_127721936_127723840)
         );
  XOR2X1 U3095 ( .A(input_times_b0_mul_componentxUMxa8_and_b2), .B(n2423), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732256_127721936_127723840)
         );
  XOR2X1 U3096 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b3), .B(n2629), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127830672_127844928_127846832)
         );
  XOR2X1 U3097 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b3), .B(n2863), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127830672_127844928_127846832)
         );
  XOR2X1 U3098 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b3), .B(n3331), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127830672_127844928_127846832)
         );
  XOR2X1 U3099 ( .A(input_times_b0_mul_componentxUMxa2_and_b3), .B(n2395), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127830672_127844928_127846832)
         );
  XOR2X1 U3100 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b4), .B(n2649), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673120_127675024_127730240)
         );
  XOR2X1 U3101 ( .A(input_times_b0_mul_componentxUMxa5_and_b4), .B(n2415), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673120_127675024_127730240)
         );
  XOR2X1 U3102 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b5), .B(n2637), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127830896_127845152_127847056)
         );
  XOR2X1 U3103 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b5), .B(n2871), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127830896_127845152_127847056)
         );
  XOR2X1 U3104 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b5), .B(n3339), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127830896_127845152_127847056)
         );
  XOR2X1 U3105 ( .A(input_times_b0_mul_componentxUMxa2_and_b5), .B(n2403), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127830896_127845152_127847056)
         );
  XOR2X1 U3106 ( .A(input_p1_times_b1_mul_componentxUMxa13_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa12_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127715536_127848576)
         );
  XOR2X1 U3107 ( .A(input_times_b0_mul_componentxUMxa13_and_b0), 
        .B(input_times_b0_mul_componentxUMxa12_and_b1), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127715536_127848576) );
  XOR2X1 U3108 ( .A(input_p2_times_b2_mul_componentxUMxa13_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa12_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127715536_127848576)
         );
  XOR2X1 U3109 ( .A(output_p2_times_a2_mul_componentxUMxa13_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa12_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127715536_127848576)
         );
  XOR2X1 U3110 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b2), .B(n2639), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127672896_127674800_127730016)
         );
  XOR2X1 U3111 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b2), .B(n2873), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127672896_127674800_127730016)
         );
  XOR2X1 U3112 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b2), .B(n3341), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127672896_127674800_127730016)
         );
  XOR2X1 U3113 ( .A(input_times_b0_mul_componentxUMxa5_and_b2), .B(n2405), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127672896_127674800_127730016)
         );
  XOR2X1 U3114 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b4), .B(n2633), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127830784_127845040_127846944)
         );
  XOR2X1 U3115 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b4), .B(n2867), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127830784_127845040_127846944)
         );
  XOR2X1 U3116 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b4), .B(n3335), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127830784_127845040_127846944)
         );
  XOR2X1 U3117 ( .A(input_times_b0_mul_componentxUMxa2_and_b4), .B(n2399), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127830784_127845040_127846944)
         );
  AND2X2 U3118 ( .A(input_p1_times_b1_mul_componentxUMxa10_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa9_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer1_127635696_127637600)
         );
  AND2X2 U3119 ( .A(input_p2_times_b2_mul_componentxUMxa10_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa9_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer1_127635696_127637600)
         );
  AND2X2 U3120 ( .A(output_p2_times_a2_mul_componentxUMxa10_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa9_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer1_127635696_127637600)
         );
  AND2X2 U3121 ( .A(input_times_b0_mul_componentxUMxa10_and_b0), 
        .B(input_times_b0_mul_componentxUMxa9_and_b1), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer1_127635696_127637600)
         );
  AND2X2 U3122 ( .A(input_p1_times_b1_mul_componentxUMxa7_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa6_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer1_127731920_127721600)
         );
  AND2X2 U3123 ( .A(input_p2_times_b2_mul_componentxUMxa7_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa6_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer1_127731920_127721600)
         );
  AND2X2 U3124 ( .A(output_p2_times_a2_mul_componentxUMxa7_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa6_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer1_127731920_127721600)
         );
  AND2X2 U3125 ( .A(input_times_b0_mul_componentxUMxa7_and_b0), 
        .B(input_times_b0_mul_componentxUMxa6_and_b1), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer1_127731920_127721600)
         );
  XOR2X1 U3126 ( .A(input_p1_times_b1_mul_componentxUMxa11_and_b0), .B(n2665), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127635808_127637712_127713408)
         );
  XOR2X1 U3127 ( .A(input_times_b0_mul_componentxUMxa11_and_b0), .B(n2431), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127635808_127637712_127713408)
         );
  XOR2X1 U3128 ( .A(input_p2_times_b2_mul_componentxUMxa11_and_b0), .B(n2899), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127635808_127637712_127713408)
         );
  XOR2X1 U3129 ( .A(output_p2_times_a2_mul_componentxUMxa11_and_b0), .B(n3367), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127635808_127637712_127713408)
         );
  XOR2X1 U3130 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b1), .B(n2635), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127672784_127674688_127729904)
         );
  XOR2X1 U3131 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b1), .B(n2869), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127672784_127674688_127729904)
         );
  XOR2X1 U3132 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b1), .B(n3337), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127672784_127674688_127729904)
         );
  XOR2X1 U3133 ( .A(input_times_b0_mul_componentxUMxa5_and_b1), .B(n2401), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127672784_127674688_127729904)
         );
  XOR2X1 U3134 ( .A(input_p1_times_b1_mul_componentxUMxa7_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa6_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127731920_127721600)
         );
  XOR2X1 U3135 ( .A(input_p2_times_b2_mul_componentxUMxa7_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa6_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127731920_127721600)
         );
  XOR2X1 U3136 ( .A(output_p2_times_a2_mul_componentxUMxa7_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa6_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127731920_127721600)
         );
  XOR2X1 U3137 ( .A(input_times_b0_mul_componentxUMxa7_and_b0), 
        .B(input_times_b0_mul_componentxUMxa6_and_b1), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127731920_127721600) );
  INVX1 U3138 ( .A(n2690), .Y(n967) );
  AOI22X1 U3139 ( .A0(input_p1_times_b1_mul_componentxUMxa10_and_b4), 
        .A1(input_p1_times_b1_mul_componentxUMxa9_and_b5), .B0(n2689), 
        .B1(input_p1_times_b1_mul_componentxUMxa11_and_b3), .Y(n2690) );
  INVX1 U3140 ( .A(n2924), .Y(n1126) );
  AOI22X1 U3141 ( .A0(input_p2_times_b2_mul_componentxUMxa10_and_b4), 
        .A1(input_p2_times_b2_mul_componentxUMxa9_and_b5), .B0(n2923), 
        .B1(input_p2_times_b2_mul_componentxUMxa11_and_b3), .Y(n2924) );
  INVX1 U3142 ( .A(n3392), .Y(n649) );
  AOI22X1 U3143 ( .A0(output_p2_times_a2_mul_componentxUMxa10_and_b4), 
        .A1(output_p2_times_a2_mul_componentxUMxa9_and_b5), .B0(n3391), 
        .B1(output_p2_times_a2_mul_componentxUMxa11_and_b3), .Y(n3392) );
  INVX1 U3144 ( .A(n2456), .Y(n808) );
  AOI22X1 U3145 ( .A0(input_times_b0_mul_componentxUMxa10_and_b4), 
        .A1(input_times_b0_mul_componentxUMxa9_and_b5), .B0(n2455), 
        .B1(input_times_b0_mul_componentxUMxa11_and_b3), .Y(n2456) );
  INVX1 U3146 ( .A(n2702), .Y(n984) );
  AOI22X1 U3147 ( .A0(input_p1_times_b1_mul_componentxUMxa13_and_b2), 
        .A1(input_p1_times_b1_mul_componentxUMxa12_and_b3), .B0(n2701), 
        .B1(input_p1_times_b1_mul_componentxUMxa14_and_b1), .Y(n2702) );
  INVX1 U3148 ( .A(n2936), .Y(n1143) );
  AOI22X1 U3149 ( .A0(input_p2_times_b2_mul_componentxUMxa13_and_b2), 
        .A1(input_p2_times_b2_mul_componentxUMxa12_and_b3), .B0(n2935), 
        .B1(input_p2_times_b2_mul_componentxUMxa14_and_b1), .Y(n2936) );
  INVX1 U3150 ( .A(n3404), .Y(n666) );
  AOI22X1 U3151 ( .A0(output_p2_times_a2_mul_componentxUMxa13_and_b2), 
        .A1(output_p2_times_a2_mul_componentxUMxa12_and_b3), .B0(n3403), 
        .B1(output_p2_times_a2_mul_componentxUMxa14_and_b1), .Y(n3404) );
  INVX1 U3152 ( .A(n2468), .Y(n825) );
  AOI22X1 U3153 ( .A0(input_times_b0_mul_componentxUMxa13_and_b2), 
        .A1(input_times_b0_mul_componentxUMxa12_and_b3), .B0(n2467), 
        .B1(input_times_b0_mul_componentxUMxa14_and_b1), .Y(n2468) );
  INVX1 U3154 ( .A(n2864), .Y(n1130) );
  AOI22X1 U3155 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b4), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b5), .B0(n2863), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b3), .Y(n2864) );
  INVX1 U3156 ( .A(n3332), .Y(n653) );
  AOI22X1 U3157 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b4), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b5), .B0(n3331), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b3), .Y(n3332) );
  INVX1 U3158 ( .A(n2642), .Y(n946) );
  AOI22X1 U3159 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b7), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b8), .B0(n2641), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b6), .Y(n2642) );
  INVX1 U3160 ( .A(n2640), .Y(n977) );
  AOI22X1 U3161 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b3), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b4), .B0(n2639), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b2), .Y(n2640) );
  INVX1 U3162 ( .A(n2870), .Y(n1142) );
  AOI22X1 U3163 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b2), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b3), .B0(n2869), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b1), .Y(n2870) );
  INVX1 U3164 ( .A(n3338), .Y(n665) );
  AOI22X1 U3165 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b2), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b3), .B0(n3337), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b1), .Y(n3338) );
  INVX1 U3166 ( .A(n2408), .Y(n787) );
  AOI22X1 U3167 ( .A0(input_times_b0_mul_componentxUMxa1_and_b7), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b8), .B0(n2407), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b6), .Y(n2408) );
  INVX1 U3168 ( .A(n2406), .Y(n818) );
  AOI22X1 U3169 ( .A0(input_times_b0_mul_componentxUMxa4_and_b3), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b4), .B0(n2405), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b2), .Y(n2406) );
  INVX1 U3170 ( .A(n2650), .Y(n963) );
  AOI22X1 U3171 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b5), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b6), .B0(n2649), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b4), .Y(n2650) );
  INVX1 U3172 ( .A(n2968), .Y(n1104) );
  AOI22X1 U3173 ( .A0(n1105), 
        .A1(input_p2_times_b2_mul_componentxUMxa9_and_b0), .B0(n2967), 
        .B1(n1128), .Y(n2968) );
  INVX1 U3174 ( .A(n2884), .Y(n1122) );
  AOI22X1 U3175 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b5), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b6), .B0(n2883), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b4), .Y(n2884) );
  INVX1 U3176 ( .A(n3436), .Y(n627) );
  AOI22X1 U3177 ( .A0(n628), 
        .A1(output_p2_times_a2_mul_componentxUMxa9_and_b0), .B0(n3435), 
        .B1(n651), .Y(n3436) );
  INVX1 U3178 ( .A(n3352), .Y(n645) );
  AOI22X1 U3179 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b5), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b6), .B0(n3351), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b4), .Y(n3352) );
  INVX1 U3180 ( .A(n2416), .Y(n804) );
  AOI22X1 U3181 ( .A0(input_times_b0_mul_componentxUMxa4_and_b5), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b6), .B0(n2415), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b4), .Y(n2416) );
  INVX1 U3182 ( .A(n2890), .Y(n1112) );
  AOI22X1 U3183 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b6), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b7), .B0(n2889), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b5), .Y(n2890) );
  INVX1 U3184 ( .A(n3358), .Y(n635) );
  AOI22X1 U3185 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b6), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b7), .B0(n3357), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b5), .Y(n3358) );
  INVX1 U3186 ( .A(n2908), .Y(n1140) );
  AOI22X1 U3187 ( .A0(input_p2_times_b2_mul_componentxUMxa10_and_b2), 
        .A1(input_p2_times_b2_mul_componentxUMxa9_and_b3), .B0(n2907), 
        .B1(input_p2_times_b2_mul_componentxUMxa11_and_b1), .Y(n2908) );
  INVX1 U3188 ( .A(n3376), .Y(n663) );
  AOI22X1 U3189 ( .A0(output_p2_times_a2_mul_componentxUMxa10_and_b2), 
        .A1(output_p2_times_a2_mul_componentxUMxa9_and_b3), .B0(n3375), 
        .B1(output_p2_times_a2_mul_componentxUMxa11_and_b1), .Y(n3376) );
  INVX1 U3190 ( .A(n2916), .Y(n1134) );
  AOI22X1 U3191 ( .A0(input_p2_times_b2_mul_componentxUMxa10_and_b3), 
        .A1(input_p2_times_b2_mul_componentxUMxa9_and_b4), .B0(n2915), 
        .B1(input_p2_times_b2_mul_componentxUMxa11_and_b2), .Y(n2916) );
  INVX1 U3192 ( .A(n3384), .Y(n657) );
  AOI22X1 U3193 ( .A0(output_p2_times_a2_mul_componentxUMxa10_and_b3), 
        .A1(output_p2_times_a2_mul_componentxUMxa9_and_b4), .B0(n3383), 
        .B1(output_p2_times_a2_mul_componentxUMxa11_and_b2), .Y(n3384) );
  INVX1 U3194 ( .A(n2746), .Y(n911) );
  AOI22X1 U3195 ( .A0(n912), 
        .A1(input_p1_times_b1_mul_componentxUMxa12_and_b0), .B0(n2745), 
        .B1(n944), .Y(n2746) );
  INVX1 U3196 ( .A(n2980), .Y(n1070) );
  AOI22X1 U3197 ( .A0(n1071), 
        .A1(input_p2_times_b2_mul_componentxUMxa12_and_b0), .B0(n2979), 
        .B1(n1103), .Y(n2980) );
  INVX1 U3198 ( .A(n3448), .Y(n593) );
  AOI22X1 U3199 ( .A0(n594), 
        .A1(output_p2_times_a2_mul_componentxUMxa12_and_b0), .B0(n3447), 
        .B1(n626), .Y(n3448) );
  INVX1 U3200 ( .A(n2512), .Y(n752) );
  AOI22X1 U3201 ( .A0(n753), .A1(input_times_b0_mul_componentxUMxa12_and_b0), 
        .B0(n2511), .B1(n785), .Y(n2512) );
  INVX1 U3202 ( .A(n2626), .Y(n985) );
  AOI22X1 U3203 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b2), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b3), .B0(n2625), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b1), .Y(n2626) );
  INVX1 U3204 ( .A(n2392), .Y(n826) );
  AOI22X1 U3205 ( .A0(input_times_b0_mul_componentxUMxa1_and_b2), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b3), .B0(n2391), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b1), .Y(n2392) );
  INVX1 U3206 ( .A(n2634), .Y(n964) );
  AOI22X1 U3207 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b5), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b6), .B0(n2633), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b4), .Y(n2634) );
  INVX1 U3208 ( .A(n2638), .Y(n956) );
  AOI22X1 U3209 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b6), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b7), .B0(n2637), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b5), .Y(n2638) );
  INVX1 U3210 ( .A(n2868), .Y(n1123) );
  AOI22X1 U3211 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b5), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b6), .B0(n2867), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b4), .Y(n2868) );
  INVX1 U3212 ( .A(n3336), .Y(n646) );
  AOI22X1 U3213 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b5), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b6), .B0(n3335), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b4), .Y(n3336) );
  INVX1 U3214 ( .A(n2400), .Y(n805) );
  AOI22X1 U3215 ( .A0(input_times_b0_mul_componentxUMxa1_and_b5), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b6), .B0(n2399), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b4), .Y(n2400) );
  INVX1 U3216 ( .A(n2404), .Y(n797) );
  AOI22X1 U3217 ( .A0(input_times_b0_mul_componentxUMxa1_and_b6), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b7), .B0(n2403), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b5), .Y(n2404) );
  INVX1 U3218 ( .A(n2880), .Y(n1148) );
  AOI22X1 U3219 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b1), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b2), .B0(n2879), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b0), .Y(n2880) );
  INVX1 U3220 ( .A(n3348), .Y(n671) );
  AOI22X1 U3221 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b1), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b2), .B0(n3347), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b0), .Y(n3348) );
  INVX1 U3222 ( .A(n2692), .Y(n991) );
  AOI22X1 U3223 ( .A0(input_p1_times_b1_mul_componentxUMxa13_and_b1), 
        .A1(input_p1_times_b1_mul_componentxUMxa12_and_b2), .B0(n2691), 
        .B1(input_p1_times_b1_mul_componentxUMxa14_and_b0), .Y(n2692) );
  INVX1 U3224 ( .A(n2926), .Y(n1150) );
  AOI22X1 U3225 ( .A0(input_p2_times_b2_mul_componentxUMxa13_and_b1), 
        .A1(input_p2_times_b2_mul_componentxUMxa12_and_b2), .B0(n2925), 
        .B1(input_p2_times_b2_mul_componentxUMxa14_and_b0), .Y(n2926) );
  INVX1 U3226 ( .A(n3394), .Y(n673) );
  AOI22X1 U3227 ( .A0(output_p2_times_a2_mul_componentxUMxa13_and_b1), 
        .A1(output_p2_times_a2_mul_componentxUMxa12_and_b2), .B0(n3393), 
        .B1(output_p2_times_a2_mul_componentxUMxa14_and_b0), .Y(n3394) );
  INVX1 U3228 ( .A(n2458), .Y(n832) );
  AOI22X1 U3229 ( .A0(input_times_b0_mul_componentxUMxa13_and_b1), 
        .A1(input_times_b0_mul_componentxUMxa12_and_b2), .B0(n2457), 
        .B1(input_times_b0_mul_componentxUMxa14_and_b0), .Y(n2458) );
  INVX1 U3230 ( .A(n2632), .Y(n990) );
  AOI22X1 U3231 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b1), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b2), .B0(n2631), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b0), .Y(n2632) );
  INVX1 U3232 ( .A(n2866), .Y(n1149) );
  AOI22X1 U3233 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b1), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b2), .B0(n2865), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b0), .Y(n2866) );
  INVX1 U3234 ( .A(n3334), .Y(n672) );
  AOI22X1 U3235 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b1), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b2), .B0(n3333), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b0), .Y(n3334) );
  INVX1 U3236 ( .A(n2398), .Y(n831) );
  AOI22X1 U3237 ( .A0(input_times_b0_mul_componentxUMxa4_and_b1), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b2), .B0(n2397), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b0), .Y(n2398) );
  INVX1 U3238 ( .A(n2644), .Y(n969) );
  AOI22X1 U3239 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b4), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b5), .B0(n2643), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b3), .Y(n2644) );
  INVX1 U3240 ( .A(n2878), .Y(n1128) );
  AOI22X1 U3241 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b4), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b5), .B0(n2877), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b3), .Y(n2878) );
  INVX1 U3242 ( .A(n3346), .Y(n651) );
  AOI22X1 U3243 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b4), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b5), .B0(n3345), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b3), .Y(n3346) );
  INVX1 U3244 ( .A(n2410), .Y(n810) );
  AOI22X1 U3245 ( .A0(input_times_b0_mul_componentxUMxa4_and_b4), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b5), .B0(n2409), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b3), .Y(n2410) );
  INVX1 U3246 ( .A(n2652), .Y(n982) );
  AOI22X1 U3247 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b2), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b3), .B0(n2651), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b1), .Y(n2652) );
  INVX1 U3248 ( .A(n2886), .Y(n1141) );
  AOI22X1 U3249 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b2), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b3), .B0(n2885), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b1), .Y(n2886) );
  INVX1 U3250 ( .A(n3354), .Y(n664) );
  AOI22X1 U3251 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b2), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b3), .B0(n3353), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b1), .Y(n3354) );
  INVX1 U3252 ( .A(n2418), .Y(n823) );
  AOI22X1 U3253 ( .A0(input_times_b0_mul_componentxUMxa7_and_b2), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b3), .B0(n2417), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b1), .Y(n2418) );
  INVX1 U3254 ( .A(n2658), .Y(n976) );
  AOI22X1 U3255 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b3), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b4), .B0(n2657), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b2), .Y(n2658) );
  INVX1 U3256 ( .A(n2892), .Y(n1135) );
  AOI22X1 U3257 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b3), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b4), .B0(n2891), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b2), .Y(n2892) );
  INVX1 U3258 ( .A(n3360), .Y(n658) );
  AOI22X1 U3259 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b3), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b4), .B0(n3359), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b2), .Y(n3360) );
  INVX1 U3260 ( .A(n2424), .Y(n817) );
  AOI22X1 U3261 ( .A0(input_times_b0_mul_componentxUMxa7_and_b3), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b4), .B0(n2423), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b2), .Y(n2424) );
  INVX1 U3262 ( .A(n2700), .Y(n961) );
  AOI22X1 U3263 ( .A0(input_p1_times_b1_mul_componentxUMxa10_and_b5), 
        .A1(input_p1_times_b1_mul_componentxUMxa9_and_b6), .B0(n2699), 
        .B1(input_p1_times_b1_mul_componentxUMxa11_and_b4), .Y(n2700) );
  INVX1 U3264 ( .A(n2466), .Y(n802) );
  AOI22X1 U3265 ( .A0(input_times_b0_mul_componentxUMxa10_and_b5), 
        .A1(input_times_b0_mul_componentxUMxa9_and_b6), .B0(n2465), 
        .B1(input_times_b0_mul_componentxUMxa11_and_b4), .Y(n2466) );
  INVX1 U3266 ( .A(n2912), .Y(n1082) );
  AOI22X1 U3267 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b9), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b10), .B0(n2911), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b8), .Y(n2912) );
  INVX1 U3268 ( .A(n3380), .Y(n605) );
  AOI22X1 U3269 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b9), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b10), .B0(n3379), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b8), .Y(n3380) );
  AOI22X1 U3270 ( .A0(input_p1_times_b1_mul_componentxUMxa13_and_b3), 
        .A1(input_p1_times_b1_mul_componentxUMxa12_and_b4), .B0(n2711), 
        .B1(input_p1_times_b1_mul_componentxUMxa14_and_b2), .Y(n2712) );
  AOI22X1 U3271 ( .A0(input_p2_times_b2_mul_componentxUMxa13_and_b3), 
        .A1(input_p2_times_b2_mul_componentxUMxa12_and_b4), .B0(n2945), 
        .B1(input_p2_times_b2_mul_componentxUMxa14_and_b2), .Y(n2946) );
  AOI22X1 U3272 ( .A0(output_p2_times_a2_mul_componentxUMxa13_and_b3), 
        .A1(output_p2_times_a2_mul_componentxUMxa12_and_b4), .B0(n3413), 
        .B1(output_p2_times_a2_mul_componentxUMxa14_and_b2), .Y(n3414) );
  AOI22X1 U3273 ( .A0(input_times_b0_mul_componentxUMxa13_and_b3), 
        .A1(input_times_b0_mul_componentxUMxa12_and_b4), .B0(n2477), 
        .B1(input_times_b0_mul_componentxUMxa14_and_b2), .Y(n2478) );
  INVX1 U3274 ( .A(n2882), .Y(n1094) );
  AOI22X1 U3275 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b8), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b9), .B0(n2881), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b7), .Y(n2882) );
  INVX1 U3276 ( .A(n2904), .Y(n1091) );
  AOI22X1 U3277 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b8), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b9), .B0(n2903), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b7), .Y(n2904) );
  INVX1 U3278 ( .A(n3350), .Y(n617) );
  AOI22X1 U3279 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b8), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b9), .B0(n3349), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b7), .Y(n3350) );
  INVX1 U3280 ( .A(n3372), .Y(n614) );
  AOI22X1 U3281 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b8), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b9), .B0(n3371), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b7), .Y(n3372) );
  INVX1 U3282 ( .A(n2922), .Y(n1102) );
  AOI22X1 U3283 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b7), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b8), .B0(n2921), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b6), .Y(n2922) );
  INVX1 U3284 ( .A(n3390), .Y(n625) );
  AOI22X1 U3285 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b7), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b8), .B0(n3389), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b6), .Y(n3390) );
  XOR2X1 U3286 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b11), .B(n2675), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831568_127845824_127847728)
         );
  XOR2X1 U3287 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b11), .B(n2909), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831568_127845824_127847728)
         );
  XOR2X1 U3288 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b11), .B(n3377), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831568_127845824_127847728)
         );
  XOR2X1 U3289 ( .A(input_times_b0_mul_componentxUMxa2_and_b11), .B(n2441), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831568_127845824_127847728)
         );
  XOR2X1 U3290 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b7), .B(n2647), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831120_127845376_127847280)
         );
  XOR2X1 U3291 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b7), .B(n2881), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831120_127845376_127847280)
         );
  XOR2X1 U3292 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b7), .B(n3349), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831120_127845376_127847280)
         );
  XOR2X1 U3293 ( .A(input_times_b0_mul_componentxUMxa2_and_b7), .B(n2413), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831120_127845376_127847280)
         );
  XOR2X1 U3294 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b9), .B(n2659), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831344_127845600_127847504)
         );
  XOR2X1 U3295 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b9), .B(n2893), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831344_127845600_127847504)
         );
  XOR2X1 U3296 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b9), .B(n3361), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831344_127845600_127847504)
         );
  XOR2X1 U3297 ( .A(input_times_b0_mul_componentxUMxa2_and_b9), .B(n2425), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831344_127845600_127847504)
         );
  XOR2X1 U3298 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b6), .B(n2921), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732704_127722384_127724288)
         );
  XOR2X1 U3299 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b6), .B(n3389), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732704_127722384_127724288)
         );
  XOR2X1 U3300 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b10), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b9), .Y(n2653) );
  XOR2X1 U3301 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b10), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b9), .Y(n2887) );
  XOR2X1 U3302 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b10), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b9), .Y(n3355) );
  XOR2X1 U3303 ( .A(input_times_b0_mul_componentxUMxa0_and_b10), 
        .B(input_times_b0_mul_componentxUMxa1_and_b9), .Y(n2419) );
  XOR2X1 U3304 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b10), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b9), .Y(n2677) );
  XOR2X1 U3305 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b10), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b9), .Y(n2911) );
  XOR2X1 U3306 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b10), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b9), .Y(n3379) );
  XOR2X1 U3307 ( .A(input_times_b0_mul_componentxUMxa3_and_b10), 
        .B(input_times_b0_mul_componentxUMxa4_and_b9), .Y(n2443) );
  XOR2X1 U3308 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b11), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b10), .Y(n2685) );
  XOR2X1 U3309 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b11), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b10), .Y(n2919) );
  XOR2X1 U3310 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b11), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b10), .Y(n3387) );
  XOR2X1 U3311 ( .A(input_times_b0_mul_componentxUMxa3_and_b11), 
        .B(input_times_b0_mul_componentxUMxa4_and_b10), .Y(n2451) );
  XOR2X1 U3312 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b11), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b10), .Y(n2659) );
  XOR2X1 U3313 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b11), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b10), .Y(n2893) );
  XOR2X1 U3314 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b11), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b10), .Y(n3361) );
  XOR2X1 U3315 ( .A(input_times_b0_mul_componentxUMxa0_and_b11), 
        .B(input_times_b0_mul_componentxUMxa1_and_b10), .Y(n2425) );
  XOR2X1 U3316 ( .A(input_p1_times_b1_mul_componentxUMxa12_and_b4), 
        .B(input_p1_times_b1_mul_componentxUMxa13_and_b3), .Y(n2711) );
  XOR2X1 U3317 ( .A(input_times_b0_mul_componentxUMxa12_and_b4), 
        .B(input_times_b0_mul_componentxUMxa13_and_b3), .Y(n2477) );
  XOR2X1 U3318 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b12), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b11), .Y(n2667) );
  XOR2X1 U3319 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b12), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b11), .Y(n2901) );
  XOR2X1 U3320 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b12), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b11), .Y(n3369) );
  XOR2X1 U3321 ( .A(input_times_b0_mul_componentxUMxa0_and_b12), 
        .B(input_times_b0_mul_componentxUMxa1_and_b11), .Y(n2433) );
  XOR2X1 U3322 ( .A(input_p2_times_b2_mul_componentxUMxa12_and_b4), 
        .B(input_p2_times_b2_mul_componentxUMxa13_and_b3), .Y(n2945) );
  XOR2X1 U3323 ( .A(output_p2_times_a2_mul_componentxUMxa12_and_b4), 
        .B(output_p2_times_a2_mul_componentxUMxa13_and_b3), .Y(n3413) );
  XOR2X1 U3324 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b13), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b12), .Y(n2675) );
  XOR2X1 U3325 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b13), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b12), .Y(n2909) );
  XOR2X1 U3326 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b13), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b12), .Y(n3377) );
  XOR2X1 U3327 ( .A(input_times_b0_mul_componentxUMxa0_and_b13), 
        .B(input_times_b0_mul_componentxUMxa1_and_b12), .Y(n2441) );
  XOR2X1 U3328 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b2), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b1), .Y(n2623) );
  XOR2X1 U3329 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b2), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b1), .Y(n2857) );
  XOR2X1 U3330 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b2), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b1), .Y(n3325) );
  XOR2X1 U3331 ( .A(input_times_b0_mul_componentxUMxa0_and_b2), 
        .B(input_times_b0_mul_componentxUMxa1_and_b1), 
        .Y(input_times_b0_mul_componentxUMxFA_127826296_127826240xn2) );
  XOR2X1 U3332 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b9), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b8), .Y(n2647) );
  XOR2X1 U3333 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b9), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b8), .Y(n2881) );
  XOR2X1 U3334 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b9), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b8), .Y(n3349) );
  XOR2X1 U3335 ( .A(input_times_b0_mul_componentxUMxa0_and_b9), 
        .B(input_times_b0_mul_componentxUMxa1_and_b8), .Y(n2413) );
  XOR2X1 U3336 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b0), .B(n992), 
        .Y(n2719) );
  XOR2X1 U3337 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b0), .B(n1151), 
        .Y(n2953) );
  XOR2X1 U3338 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b0), .B(n674), 
        .Y(n3421) );
  XOR2X1 U3339 ( .A(input_times_b0_mul_componentxUMxa3_and_b0), .B(n833), 
        .Y(n2485) );
  XOR2X1 U3340 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b9), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b8), .Y(n2669) );
  XOR2X1 U3341 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b9), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b8), .Y(n2903) );
  XOR2X1 U3342 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b9), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b8), .Y(n3371) );
  XOR2X1 U3343 ( .A(input_times_b0_mul_componentxUMxa3_and_b9), 
        .B(input_times_b0_mul_componentxUMxa4_and_b8), .Y(n2435) );
  XOR2X1 U3344 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b8), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b7), .Y(n2661) );
  XOR2X1 U3345 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b8), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b7), .Y(n2895) );
  XOR2X1 U3346 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b8), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b7), .Y(n3363) );
  XOR2X1 U3347 ( .A(input_times_b0_mul_componentxUMxa3_and_b8), 
        .B(input_times_b0_mul_componentxUMxa4_and_b7), .Y(n2427) );
  XOR2X1 U3348 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b7), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b6), .Y(n2679) );
  XOR2X1 U3349 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b7), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b6), .Y(n2913) );
  XOR2X1 U3350 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b7), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b6), .Y(n3381) );
  XOR2X1 U3351 ( .A(input_times_b0_mul_componentxUMxa6_and_b7), 
        .B(input_times_b0_mul_componentxUMxa7_and_b6), .Y(n2445) );
  XOR2X1 U3352 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b8), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b7), .Y(n2921) );
  XOR2X1 U3353 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b8), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b7), .Y(n3389) );
  XOR2X1 U3354 ( .A(input_p1_times_b1_mul_componentxUMxa9_and_b6), 
        .B(input_p1_times_b1_mul_componentxUMxa10_and_b5), .Y(n2699) );
  XOR2X1 U3355 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b9), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b8), .Y(n2697) );
  XOR2X1 U3356 ( .A(input_p2_times_b2_mul_componentxUMxa9_and_b6), 
        .B(input_p2_times_b2_mul_componentxUMxa10_and_b5), .Y(n2933) );
  XOR2X1 U3357 ( .A(output_p2_times_a2_mul_componentxUMxa9_and_b6), 
        .B(output_p2_times_a2_mul_componentxUMxa10_and_b5), .Y(n3401) );
  XOR2X1 U3358 ( .A(input_times_b0_mul_componentxUMxa9_and_b6), 
        .B(input_times_b0_mul_componentxUMxa10_and_b5), .Y(n2465) );
  XOR2X1 U3359 ( .A(input_times_b0_mul_componentxUMxa6_and_b9), 
        .B(input_times_b0_mul_componentxUMxa7_and_b8), .Y(n2463) );
  XOR2X1 U3360 ( .A(input_p1_times_b1_mul_componentxUMxa9_and_b7), 
        .B(input_p1_times_b1_mul_componentxUMxa10_and_b6), .Y(n2709) );
  XOR2X1 U3361 ( .A(input_p2_times_b2_mul_componentxUMxa9_and_b7), 
        .B(input_p2_times_b2_mul_componentxUMxa10_and_b6), .Y(n2943) );
  XOR2X1 U3362 ( .A(output_p2_times_a2_mul_componentxUMxa9_and_b7), 
        .B(output_p2_times_a2_mul_componentxUMxa10_and_b6), .Y(n3411) );
  XOR2X1 U3363 ( .A(input_times_b0_mul_componentxUMxa9_and_b7), 
        .B(input_times_b0_mul_componentxUMxa10_and_b6), .Y(n2475) );
  XOR2X1 U3364 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b0), .B(n2631), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127672672_127674576_127729792)
         );
  XOR2X1 U3365 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b0), .B(n2865), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127672672_127674576_127729792)
         );
  XOR2X1 U3366 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b0), .B(n3333), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127672672_127674576_127729792)
         );
  XOR2X1 U3367 ( .A(input_times_b0_mul_componentxUMxa5_and_b0), .B(n2397), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127672672_127674576_127729792)
         );
  XOR2X1 U3368 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b5), .B(n2679), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732592_127722272_127724176)
         );
  XOR2X1 U3369 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b5), .B(n2913), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732592_127722272_127724176)
         );
  XOR2X1 U3370 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b5), .B(n3381), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732592_127722272_127724176)
         );
  XOR2X1 U3371 ( .A(input_times_b0_mul_componentxUMxa8_and_b5), .B(n2445), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732592_127722272_127724176)
         );
  XOR2X1 U3372 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b8), .B(n2653), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831232_127845488_127847392)
         );
  XOR2X1 U3373 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b8), .B(n2887), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831232_127845488_127847392)
         );
  XOR2X1 U3374 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b8), .B(n3355), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831232_127845488_127847392)
         );
  XOR2X1 U3375 ( .A(input_times_b0_mul_componentxUMxa2_and_b8), .B(n2419), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831232_127845488_127847392)
         );
  XOR2X1 U3376 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b7), .B(n2669), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673456_127675360_127730576)
         );
  XOR2X1 U3377 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b7), .B(n2903), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673456_127675360_127730576)
         );
  XOR2X1 U3378 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b7), .B(n3371), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673456_127675360_127730576)
         );
  XOR2X1 U3379 ( .A(input_times_b0_mul_componentxUMxa5_and_b7), .B(n2435), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673456_127675360_127730576)
         );
  XOR2X1 U3380 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b9), .B(n2685), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673680_127675584_127730800)
         );
  XOR2X1 U3381 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b9), .B(n2919), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673680_127675584_127730800)
         );
  XOR2X1 U3382 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b9), .B(n3387), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673680_127675584_127730800)
         );
  XOR2X1 U3383 ( .A(input_times_b0_mul_componentxUMxa5_and_b9), .B(n2451), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673680_127675584_127730800)
         );
  XOR2X1 U3384 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b10), .B(n2667), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831456_127845712_127847616)
         );
  XOR2X1 U3385 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b10), .B(n2901), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831456_127845712_127847616)
         );
  XOR2X1 U3386 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b10), .B(n3369), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831456_127845712_127847616)
         );
  XOR2X1 U3387 ( .A(input_times_b0_mul_componentxUMxa2_and_b10), .B(n2433), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831456_127845712_127847616)
         );
  XOR2X1 U3388 ( .A(input_p1_times_b1_mul_componentxUMxa11_and_b5), .B(n2709), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127636368_127638272_127713968)
         );
  XOR2X1 U3389 ( .A(input_times_b0_mul_componentxUMxa11_and_b5), .B(n2475), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127636368_127638272_127713968)
         );
  XOR2X1 U3390 ( .A(input_p2_times_b2_mul_componentxUMxa11_and_b5), .B(n2943), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127636368_127638272_127713968)
         );
  XOR2X1 U3391 ( .A(output_p2_times_a2_mul_componentxUMxa11_and_b5), .B(n3411), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127636368_127638272_127713968)
         );
  OAI2BB2X1 U3392 ( .B0(n133), .B1(n1260), .A0N(output_previous_2[17]), 
        .A1N(n319), .Y(n4672) );
  XOR2X1 U3393 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b1), .B(n2625), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127830448_127844704_127846608)
         );
  XOR2X1 U3394 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b1), .B(n2859), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127830448_127844704_127846608)
         );
  XOR2X1 U3395 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b1), .B(n3327), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127830448_127844704_127846608)
         );
  XOR2X1 U3396 ( .A(input_times_b0_mul_componentxUMxa2_and_b1), .B(n2391), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127830448_127844704_127846608)
         );
  XOR2X1 U3397 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b4), .B(n2883), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673120_127675024_127730240)
         );
  XOR2X1 U3398 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b4), .B(n3351), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673120_127675024_127730240)
         );
  XOR2X1 U3399 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b6), .B(n2661), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673344_127675248_127730464)
         );
  XOR2X1 U3400 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b6), .B(n2895), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673344_127675248_127730464)
         );
  XOR2X1 U3401 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b6), .B(n3363), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673344_127675248_127730464)
         );
  XOR2X1 U3402 ( .A(input_times_b0_mul_componentxUMxa5_and_b6), .B(n2427), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673344_127675248_127730464)
         );
  XOR2X1 U3403 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b7), .B(n2697), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732816_127722496_127724400)
         );
  XOR2X1 U3404 ( .A(input_times_b0_mul_componentxUMxa8_and_b7), .B(n2463), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732816_127722496_127724400)
         );
  XOR2X1 U3405 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b8), .B(n2677), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673568_127675472_127730688)
         );
  XOR2X1 U3406 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b8), .B(n2911), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673568_127675472_127730688)
         );
  XOR2X1 U3407 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b8), .B(n3379), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673568_127675472_127730688)
         );
  XOR2X1 U3408 ( .A(input_times_b0_mul_componentxUMxa5_and_b8), .B(n2443), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673568_127675472_127730688)
         );
  XOR2X1 U3409 ( .A(input_p1_times_b1_mul_componentxUMxa4_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa3_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127672560_127674464)
         );
  XOR2X1 U3410 ( .A(input_p2_times_b2_mul_componentxUMxa4_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa3_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127672560_127674464)
         );
  XOR2X1 U3411 ( .A(output_p2_times_a2_mul_componentxUMxa4_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa3_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127672560_127674464)
         );
  XOR2X1 U3412 ( .A(input_times_b0_mul_componentxUMxa4_and_b0), 
        .B(input_times_b0_mul_componentxUMxa3_and_b1), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127672560_127674464) );
  XOR2X1 U3413 ( .A(input_p1_times_b1_mul_componentxUMxa11_and_b4), .B(n2699), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127636256_127638160_127713856)
         );
  XOR2X1 U3414 ( .A(input_times_b0_mul_componentxUMxa11_and_b4), .B(n2465), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127636256_127638160_127713856)
         );
  XOR2X1 U3415 ( .A(input_p2_times_b2_mul_componentxUMxa11_and_b4), .B(n2933), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127636256_127638160_127713856)
         );
  XOR2X1 U3416 ( .A(output_p2_times_a2_mul_componentxUMxa11_and_b4), .B(n3401), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127636256_127638160_127713856)
         );
  XOR2X1 U3417 ( .A(input_p1_times_b1_mul_componentxUMxa14_and_b2), .B(n2711), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127715872_127848912_127850816)
         );
  XOR2X1 U3418 ( .A(input_times_b0_mul_componentxUMxa14_and_b2), .B(n2477), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127715872_127848912_127850816)
         );
  XOR2X1 U3419 ( .A(input_p2_times_b2_mul_componentxUMxa14_and_b2), .B(n2945), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127715872_127848912_127850816)
         );
  XOR2X1 U3420 ( .A(output_p2_times_a2_mul_componentxUMxa14_and_b2), .B(n3413), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127715872_127848912_127850816)
         );
  XOR2X1 U3421 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b3), .B(n2663), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732368_127722048_127723952)
         );
  XOR2X1 U3422 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b3), .B(n2897), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732368_127722048_127723952)
         );
  XOR2X1 U3423 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b3), .B(n3365), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732368_127722048_127723952)
         );
  XOR2X1 U3424 ( .A(input_times_b0_mul_componentxUMxa8_and_b3), .B(n2429), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732368_127722048_127723952)
         );
  XOR2X1 U3425 ( .A(input_p1_times_b1_mul_componentxUMxa14_and_b1), .B(n2701), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127715760_127848800_127850704)
         );
  XOR2X1 U3426 ( .A(input_times_b0_mul_componentxUMxa14_and_b1), .B(n2467), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127715760_127848800_127850704)
         );
  XOR2X1 U3427 ( .A(input_p2_times_b2_mul_componentxUMxa14_and_b1), .B(n2935), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127715760_127848800_127850704)
         );
  XOR2X1 U3428 ( .A(output_p2_times_a2_mul_componentxUMxa14_and_b1), .B(n3403), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127715760_127848800_127850704)
         );
  XOR2X1 U3429 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b0), .B(n2623), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127830336_127844592_127846496)
         );
  XOR2X1 U3430 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b0), .B(n2857), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127830336_127844592_127846496)
         );
  XOR2X1 U3431 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b0), .B(n3325), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127830336_127844592_127846496)
         );
  XOR2X1 U3432 ( .A(input_times_b0_mul_componentxUMxa2_and_b0), 
        .B(input_times_b0_mul_componentxUMxFA_127826296_127826240xn2), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127830336_127844592_127846496)
         );
  XOR2X1 U3433 ( .A(input_p1_times_b1_mul_componentxUMxa16_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa15_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127627504_127629408)
         );
  XOR2X1 U3434 ( .A(input_times_b0_mul_componentxUMxa16_and_b0), 
        .B(input_times_b0_mul_componentxUMxa15_and_b1), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127627504_127629408) );
  XOR2X1 U3435 ( .A(input_p2_times_b2_mul_componentxUMxa16_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa15_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127627504_127629408)
         );
  XOR2X1 U3436 ( .A(output_p2_times_a2_mul_componentxUMxa16_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa15_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127627504_127629408)
         );
  XOR2X1 U3437 ( .A(n2710), .B(n2712), .Y(n2776) );
  AOI22X1 U3438 ( .A0(input_p1_times_b1_mul_componentxUMxa10_and_b6), 
        .A1(input_p1_times_b1_mul_componentxUMxa9_and_b7), .B0(n2709), 
        .B1(input_p1_times_b1_mul_componentxUMxa11_and_b5), .Y(n2710) );
  XOR2X1 U3439 ( .A(n2944), .B(n2946), .Y(n3010) );
  AOI22X1 U3440 ( .A0(input_p2_times_b2_mul_componentxUMxa10_and_b6), 
        .A1(input_p2_times_b2_mul_componentxUMxa9_and_b7), .B0(n2943), 
        .B1(input_p2_times_b2_mul_componentxUMxa11_and_b5), .Y(n2944) );
  XOR2X1 U3441 ( .A(n3412), .B(n3414), .Y(n3478) );
  AOI22X1 U3442 ( .A0(output_p2_times_a2_mul_componentxUMxa10_and_b6), 
        .A1(output_p2_times_a2_mul_componentxUMxa9_and_b7), .B0(n3411), 
        .B1(output_p2_times_a2_mul_componentxUMxa11_and_b5), .Y(n3412) );
  XOR2X1 U3443 ( .A(n2476), .B(n2478), .Y(n2542) );
  AOI22X1 U3444 ( .A0(input_times_b0_mul_componentxUMxa10_and_b6), 
        .A1(input_times_b0_mul_componentxUMxa9_and_b7), .B0(n2475), 
        .B1(input_times_b0_mul_componentxUMxa11_and_b5), .Y(n2476) );
  INVX1 U3445 ( .A(n2660), .Y(n912) );
  AOI22X1 U3446 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b10), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b11), .B0(n2659), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b9), .Y(n2660) );
  INVX1 U3447 ( .A(n2894), .Y(n1071) );
  AOI22X1 U3448 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b10), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b11), .B0(n2893), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b9), .Y(n2894) );
  INVX1 U3449 ( .A(n3362), .Y(n594) );
  AOI22X1 U3450 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b10), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b11), .B0(n3361), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b9), .Y(n3362) );
  INVX1 U3451 ( .A(n2426), .Y(n753) );
  AOI22X1 U3452 ( .A0(input_times_b0_mul_componentxUMxa1_and_b10), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b11), .B0(n2425), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b9), .Y(n2426) );
  INVX1 U3453 ( .A(n2678), .Y(n923) );
  AOI22X1 U3454 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b9), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b10), .B0(n2677), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b8), .Y(n2678) );
  INVX1 U3455 ( .A(n2444), .Y(n764) );
  AOI22X1 U3456 ( .A0(input_times_b0_mul_componentxUMxa4_and_b9), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b10), .B0(n2443), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b8), .Y(n2444) );
  INVX1 U3457 ( .A(n2876), .Y(n1105) );
  AOI22X1 U3458 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b7), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b8), .B0(n2875), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b6), .Y(n2876) );
  INVX1 U3459 ( .A(n3344), .Y(n628) );
  AOI22X1 U3460 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b7), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b8), .B0(n3343), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b6), .Y(n3344) );
  INVX1 U3461 ( .A(n2624), .Y(n992) );
  AOI22X1 U3462 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b1), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b2), .B0(n2623), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b0), .Y(n2624) );
  INVX1 U3463 ( .A(n2858), .Y(n1151) );
  AOI22X1 U3464 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b1), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b2), .B0(n2857), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b0), .Y(n2858) );
  INVX1 U3465 ( .A(n3326), .Y(n674) );
  AOI22X1 U3466 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b1), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b2), .B0(n3325), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b0), .Y(n3326) );
  INVX1 U3467 ( .A(input_times_b0_mul_componentxUMxFA_127826296_127826240xn3), 
        .Y(n833) );
  AOI22X1 U3468 ( .A0(input_times_b0_mul_componentxUMxa1_and_b1), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b2), 
        .B0(input_times_b0_mul_componentxUMxFA_127826296_127826240xn2), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b0), 
        .Y(input_times_b0_mul_componentxUMxFA_127826296_127826240xn3) );
  INVX1 U3469 ( .A(n2670), .Y(n932) );
  AOI22X1 U3470 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b8), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b9), .B0(n2669), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b7), .Y(n2670) );
  INVX1 U3471 ( .A(n2436), .Y(n773) );
  AOI22X1 U3472 ( .A0(input_times_b0_mul_componentxUMxa4_and_b8), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b9), .B0(n2435), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b7), .Y(n2436) );
  INVX1 U3473 ( .A(n2654), .Y(n927) );
  AOI22X1 U3474 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b9), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b10), .B0(n2653), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b8), .Y(n2654) );
  INVX1 U3475 ( .A(n2888), .Y(n1086) );
  AOI22X1 U3476 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b9), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b10), .B0(n2887), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b8), .Y(n2888) );
  INVX1 U3477 ( .A(n3356), .Y(n609) );
  AOI22X1 U3478 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b9), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b10), .B0(n3355), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b8), .Y(n3356) );
  INVX1 U3479 ( .A(n2420), .Y(n768) );
  AOI22X1 U3480 ( .A0(input_times_b0_mul_componentxUMxa1_and_b9), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b10), .B0(n2419), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b8), .Y(n2420) );
  INVX1 U3481 ( .A(n2668), .Y(n904) );
  AOI22X1 U3482 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b11), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b12), .B0(n2667), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b10), .Y(n2668) );
  INVX1 U3483 ( .A(n2902), .Y(n1063) );
  AOI22X1 U3484 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b11), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b12), .B0(n2901), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b10), .Y(n2902) );
  INVX1 U3485 ( .A(n3370), .Y(n586) );
  AOI22X1 U3486 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b11), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b12), .B0(n3369), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b10), .Y(n3370) );
  INVX1 U3487 ( .A(n2434), .Y(n745) );
  AOI22X1 U3488 ( .A0(input_times_b0_mul_componentxUMxa1_and_b11), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b12), .B0(n2433), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b10), .Y(n2434) );
  INVX1 U3489 ( .A(n2934), .Y(n1120) );
  AOI22X1 U3490 ( .A0(input_p2_times_b2_mul_componentxUMxa10_and_b5), 
        .A1(input_p2_times_b2_mul_componentxUMxa9_and_b6), .B0(n2933), 
        .B1(input_p2_times_b2_mul_componentxUMxa11_and_b4), .Y(n2934) );
  INVX1 U3491 ( .A(n3402), .Y(n643) );
  AOI22X1 U3492 ( .A0(output_p2_times_a2_mul_componentxUMxa10_and_b5), 
        .A1(output_p2_times_a2_mul_componentxUMxa9_and_b6), .B0(n3401), 
        .B1(output_p2_times_a2_mul_componentxUMxa11_and_b4), .Y(n3402) );
  INVX1 U3493 ( .A(n2676), .Y(n902) );
  AOI22X1 U3494 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b12), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b13), .B0(n2675), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b11), .Y(n2676) );
  INVX1 U3495 ( .A(n2910), .Y(n1061) );
  AOI22X1 U3496 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b12), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b13), .B0(n2909), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b11), .Y(n2910) );
  INVX1 U3497 ( .A(n3378), .Y(n584) );
  AOI22X1 U3498 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b12), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b13), .B0(n3377), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b11), .Y(n3378) );
  INVX1 U3499 ( .A(n2442), .Y(n743) );
  AOI22X1 U3500 ( .A0(input_times_b0_mul_componentxUMxa1_and_b12), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b13), .B0(n2441), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b11), .Y(n2442) );
  XOR2X1 U3501 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127627616_127629520_127824000), 
        .B(n2778), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128199816_128200040_128199984)
         );
  XOR2X1 U3502 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127636480_127638384_127714080), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127715984_127849024_127850928), 
        .Y(n2778) );
  XOR2X1 U3503 ( .A(input_p1_times_b1_mul_componentxUMxa17_and_b0), .B(n2718), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127627616_127629520_127824000)
         );
  XOR2X1 U3504 ( .A(input_p1_times_b1_mul_componentxUMxa11_and_b6), .B(n2716), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127636480_127638384_127714080)
         );
  XOR2X1 U3505 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127627616_127629520_127824000), 
        .B(n3012), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128199816_128200040_128199984)
         );
  XOR2X1 U3506 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127636480_127638384_127714080), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127715984_127849024_127850928), 
        .Y(n3012) );
  XOR2X1 U3507 ( .A(input_p2_times_b2_mul_componentxUMxa17_and_b0), .B(n2952), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127627616_127629520_127824000)
         );
  XOR2X1 U3508 ( .A(input_p2_times_b2_mul_componentxUMxa11_and_b6), .B(n2950), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127636480_127638384_127714080)
         );
  XOR2X1 U3509 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127627616_127629520_127824000), 
        .B(n3480), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128199816_128200040_128199984)
         );
  XOR2X1 U3510 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127636480_127638384_127714080), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127715984_127849024_127850928), 
        .Y(n3480) );
  XOR2X1 U3511 ( .A(output_p2_times_a2_mul_componentxUMxa17_and_b0), .B(n3420), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127627616_127629520_127824000)
         );
  XOR2X1 U3512 ( .A(output_p2_times_a2_mul_componentxUMxa11_and_b6), .B(n3418), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127636480_127638384_127714080)
         );
  XOR2X1 U3513 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127627616_127629520_127824000), 
        .B(n2544), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128199816_128200040_128199984)
         );
  XOR2X1 U3514 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127636480_127638384_127714080), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127715984_127849024_127850928), 
        .Y(n2544) );
  XOR2X1 U3515 ( .A(input_times_b0_mul_componentxUMxa17_and_b0), .B(n2484), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127627616_127629520_127824000)
         );
  XOR2X1 U3516 ( .A(input_times_b0_mul_componentxUMxa11_and_b6), .B(n2482), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127636480_127638384_127714080)
         );
  INVX1 U3517 ( .A(n2648), .Y(n935) );
  AOI22X1 U3518 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b8), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b9), .B0(n2647), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b7), .Y(n2648) );
  INVX1 U3519 ( .A(n2414), .Y(n776) );
  AOI22X1 U3520 ( .A0(input_times_b0_mul_componentxUMxa1_and_b8), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b9), .B0(n2413), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b7), .Y(n2414) );
  INVX1 U3521 ( .A(n2688), .Y(n943) );
  AOI22X1 U3522 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b7), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b8), .B0(n2687), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b6), .Y(n2688) );
  INVX1 U3523 ( .A(n2454), .Y(n784) );
  AOI22X1 U3524 ( .A0(input_times_b0_mul_componentxUMxa7_and_b7), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b8), .B0(n2453), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b6), .Y(n2454) );
  INVX1 U3525 ( .A(n2764), .Y(n886) );
  AOI22X1 U3526 ( .A0(n919), 
        .A1(input_p1_times_b1_mul_componentxUMxa15_and_b0), .B0(n2763), 
        .B1(n887), .Y(n2764) );
  INVX1 U3527 ( .A(n2998), .Y(n1045) );
  AOI22X1 U3528 ( .A0(n1078), 
        .A1(input_p2_times_b2_mul_componentxUMxa15_and_b0), .B0(n2997), 
        .B1(n1046), .Y(n2998) );
  INVX1 U3529 ( .A(n3466), .Y(n568) );
  AOI22X1 U3530 ( .A0(n601), 
        .A1(output_p2_times_a2_mul_componentxUMxa15_and_b0), .B0(n3465), 
        .B1(n569), .Y(n3466) );
  INVX1 U3531 ( .A(n2530), .Y(n727) );
  AOI22X1 U3532 ( .A0(n760), .A1(input_times_b0_mul_componentxUMxa15_and_b0), 
        .B0(n2529), .B1(n728), .Y(n2530) );
  INVX1 U3533 ( .A(n2662), .Y(n944) );
  AOI22X1 U3534 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b7), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b8), .B0(n2661), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b6), .Y(n2662) );
  INVX1 U3535 ( .A(n2672), .Y(n962) );
  AOI22X1 U3536 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b5), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b6), .B0(n2671), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b4), .Y(n2672) );
  INVX1 U3537 ( .A(n2896), .Y(n1103) );
  AOI22X1 U3538 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b7), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b8), .B0(n2895), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b6), .Y(n2896) );
  INVX1 U3539 ( .A(n2906), .Y(n1121) );
  AOI22X1 U3540 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b5), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b6), .B0(n2905), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b4), .Y(n2906) );
  INVX1 U3541 ( .A(n3364), .Y(n626) );
  AOI22X1 U3542 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b7), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b8), .B0(n3363), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b6), .Y(n3364) );
  INVX1 U3543 ( .A(n3374), .Y(n644) );
  AOI22X1 U3544 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b5), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b6), .B0(n3373), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b4), .Y(n3374) );
  INVX1 U3545 ( .A(n2428), .Y(n785) );
  AOI22X1 U3546 ( .A0(input_times_b0_mul_componentxUMxa4_and_b7), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b8), .B0(n2427), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b6), .Y(n2428) );
  INVX1 U3547 ( .A(n2438), .Y(n803) );
  AOI22X1 U3548 ( .A0(input_times_b0_mul_componentxUMxa7_and_b5), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b6), .B0(n2437), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b4), .Y(n2438) );
  INVX1 U3549 ( .A(n2680), .Y(n951) );
  AOI22X1 U3550 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b6), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b7), .B0(n2679), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b5), .Y(n2680) );
  INVX1 U3551 ( .A(n2914), .Y(n1110) );
  AOI22X1 U3552 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b6), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b7), .B0(n2913), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b5), .Y(n2914) );
  INVX1 U3553 ( .A(n3382), .Y(n633) );
  AOI22X1 U3554 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b6), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b7), .B0(n3381), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b5), .Y(n3382) );
  INVX1 U3555 ( .A(n2446), .Y(n792) );
  AOI22X1 U3556 ( .A0(input_times_b0_mul_componentxUMxa7_and_b6), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b7), .B0(n2445), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b5), .Y(n2446) );
  INVX1 U3557 ( .A(n2720), .Y(n987) );
  AOI22X1 U3558 ( .A0(n992), .A1(input_p1_times_b1_mul_componentxUMxa3_and_b0), 
        .B0(n2719), 
        .B1(input_p1_times_b1_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .Y(n2720) );
  INVX1 U3559 ( .A(n2954), .Y(n1146) );
  AOI22X1 U3560 ( .A0(n1151), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b0), .B0(n2953), 
        .B1(input_p2_times_b2_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .Y(n2954) );
  INVX1 U3561 ( .A(n3422), .Y(n669) );
  AOI22X1 U3562 ( .A0(n674), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b0), .B0(n3421), 
        .B1(output_p2_times_a2_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .Y(n3422) );
  INVX1 U3563 ( .A(n2486), .Y(n828) );
  AOI22X1 U3564 ( .A0(n833), .A1(input_times_b0_mul_componentxUMxa3_and_b0), 
        .B0(n2485), 
        .B1(input_times_b0_mul_componentxUMxsum_layer1_127830448_127844704_127846608), 
        .Y(n2486) );
  AND2X2 U3565 ( .A(input_p1_times_b1_mul_componentxUMxa16_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa15_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer1_127627504_127629408)
         );
  AND2X2 U3566 ( .A(input_times_b0_mul_componentxUMxa16_and_b0), 
        .B(input_times_b0_mul_componentxUMxa15_and_b1), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer1_127627504_127629408)
         );
  AND2X2 U3567 ( .A(input_p2_times_b2_mul_componentxUMxa16_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa15_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer1_127627504_127629408)
         );
  AND2X2 U3568 ( .A(output_p2_times_a2_mul_componentxUMxa16_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa15_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer1_127627504_127629408)
         );
  INVX1 U3569 ( .A(n2696), .Y(n879) );
  AOI22X1 U3570 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b11), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b12), .B0(n2695), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b10), .Y(n2696) );
  INVX1 U3571 ( .A(n2462), .Y(n720) );
  AOI22X1 U3572 ( .A0(input_times_b0_mul_componentxUMxa4_and_b11), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b12), .B0(n2461), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b10), .Y(n2462) );
  INVX1 U3573 ( .A(n2708), .Y(n922) );
  AOI22X1 U3574 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b9), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b10), .B0(n2707), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b8), .Y(n2708) );
  INVX1 U3575 ( .A(n2474), .Y(n763) );
  AOI22X1 U3576 ( .A0(input_times_b0_mul_componentxUMxa7_and_b9), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b10), .B0(n2473), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b8), .Y(n2474) );
  INVX1 U3577 ( .A(n4449), .Y(n993) );
  AOI22XL U3578 ( .A0(input_p1_times_b1_mul_componentxUMxfirst_vector[2]), 
        .A1(n125), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[2]), 
        .B1(n4442), .Y(n4449) );
  XNOR2X1 U3579 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[2]), 
        .B(n3718), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[2]) );
  NOR2X1 U3580 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[0]), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[1]), .Y(n3718) );
  INVX1 U3581 ( .A(n4502), .Y(n1152) );
  AOI22XL U3582 ( .A0(input_p2_times_b2_mul_componentxUMxfirst_vector[2]), 
        .A1(n129), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[2]), 
        .B1(n4495), .Y(n4502) );
  XNOR2X1 U3583 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[2]), 
        .B(n3766), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[2]) );
  NOR2X1 U3584 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[0]), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[1]), .Y(n3766) );
  INVX1 U3585 ( .A(n4608), .Y(n675) );
  AOI22XL U3586 ( .A0(output_p2_times_a2_mul_componentxUMxfirst_vector[2]), 
        .A1(n117), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[2]), 
        .B1(n4601), .Y(n4608) );
  XNOR2X1 U3587 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[2]), 
        .B(n3862), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[2]) );
  NOR2X1 U3588 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[0]), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[1]), .Y(n3862) );
  INVX1 U3589 ( .A(input_times_b0_mul_componentxn98), .Y(n834) );
  AOI22XL U3590 ( .A0(input_times_b0_mul_componentxUMxfirst_vector[2]), 
        .A1(n121), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[2]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn98) );
  XNOR2X1 U3591 ( .A(input_times_b0_mul_componentxUMxfirst_vector[2]), 
        .B(n3670), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[2]) );
  NOR2X1 U3592 ( .A(input_times_b0_mul_componentxUMxfirst_vector[0]), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[1]), .Y(n3670) );
  XOR2X1 U3593 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b10), .B(n2695), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673792_127675696_127730912)
         );
  XOR2X1 U3594 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b10), .B(n2929), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673792_127675696_127730912)
         );
  XOR2X1 U3595 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b10), .B(n3397), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673792_127675696_127730912)
         );
  XOR2X1 U3596 ( .A(input_times_b0_mul_componentxUMxa5_and_b10), .B(n2461), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673792_127675696_127730912)
         );
  XOR2X1 U3597 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b8), .B(n2707), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127732928_127722608_127724512)
         );
  XOR2X1 U3598 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b8), .B(n2941), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732928_127722608_127724512)
         );
  XOR2X1 U3599 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b8), .B(n3409), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732928_127722608_127724512)
         );
  XOR2X1 U3600 ( .A(input_times_b0_mul_componentxUMxa8_and_b8), .B(n2473), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127732928_127722608_127724512)
         );
  XOR2X1 U3601 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b10), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b9), .Y(n2707) );
  XOR2X1 U3602 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b10), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b9), .Y(n2941) );
  XOR2X1 U3603 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b10), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b9), .Y(n3409) );
  XOR2X1 U3604 ( .A(input_times_b0_mul_componentxUMxa6_and_b10), 
        .B(input_times_b0_mul_componentxUMxa7_and_b9), .Y(n2473) );
  XOR2X1 U3605 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b12), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b11), .Y(n2695) );
  XOR2X1 U3606 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b12), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b11), .Y(n2929) );
  XOR2X1 U3607 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b12), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b11), .Y(n3397) );
  XOR2X1 U3608 ( .A(input_times_b0_mul_componentxUMxa3_and_b12), 
        .B(input_times_b0_mul_componentxUMxa4_and_b11), .Y(n2461) );
  XOR2X1 U3609 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b13), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b12), .Y(n2705) );
  XOR2X1 U3610 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b13), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b12), .Y(n2939) );
  XOR2X1 U3611 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b13), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b12), .Y(n3407) );
  XOR2X1 U3612 ( .A(input_times_b0_mul_componentxUMxa3_and_b13), 
        .B(input_times_b0_mul_componentxUMxa4_and_b12), .Y(n2471) );
  XOR2X1 U3613 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b14), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b13), .Y(n2683) );
  XOR2X1 U3614 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b14), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b13), .Y(n2917) );
  XOR2X1 U3615 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b14), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b13), .Y(n3385) );
  XOR2X1 U3616 ( .A(input_times_b0_mul_componentxUMxa0_and_b14), 
        .B(input_times_b0_mul_componentxUMxa1_and_b13), .Y(n2449) );
  XOR2X1 U3617 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b15), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b14), .Y(n2693) );
  XOR2X1 U3618 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b15), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b14), .Y(n2927) );
  XOR2X1 U3619 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b15), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b14), .Y(n3395) );
  XOR2X1 U3620 ( .A(input_times_b0_mul_componentxUMxa0_and_b15), 
        .B(input_times_b0_mul_componentxUMxa1_and_b14), .Y(n2459) );
  XOR2X1 U3621 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b16), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b15), .Y(n2703) );
  XOR2X1 U3622 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b16), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b15), .Y(n2937) );
  XOR2X1 U3623 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b16), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b15), .Y(n3405) );
  XOR2X1 U3624 ( .A(input_times_b0_mul_componentxUMxa0_and_b16), 
        .B(input_times_b0_mul_componentxUMxa1_and_b15), .Y(n2469) );
  XOR2X1 U3625 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b9), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b8), .Y(n2931) );
  XOR2X1 U3626 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b9), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b8), .Y(n3399) );
  OR3XL U3627 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[1]), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[2]), 
        .C(input_p1_times_b1_mul_componentxUMxfirst_vector[0]), .Y(n3717) );
  OR3XL U3628 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[1]), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[2]), 
        .C(input_p2_times_b2_mul_componentxUMxfirst_vector[0]), .Y(n3765) );
  OR3XL U3629 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[1]), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[2]), 
        .C(output_p2_times_a2_mul_componentxUMxfirst_vector[0]), .Y(n3861) );
  OR3XL U3630 ( .A(input_times_b0_mul_componentxUMxfirst_vector[1]), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[2]), 
        .C(input_times_b0_mul_componentxUMxfirst_vector[0]), .Y(n3669) );
  XOR2X1 U3631 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b11), .B(n2705), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127673904_127675808_127731024)
         );
  XOR2X1 U3632 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b11), .B(n2939), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127673904_127675808_127731024)
         );
  XOR2X1 U3633 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b11), .B(n3407), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127673904_127675808_127731024)
         );
  XOR2X1 U3634 ( .A(input_times_b0_mul_componentxUMxa5_and_b11), .B(n2471), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127673904_127675808_127731024)
         );
  XOR2X1 U3635 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b13), .B(n2693), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831792_127846048_127847952)
         );
  XOR2X1 U3636 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b13), .B(n2927), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831792_127846048_127847952)
         );
  XOR2X1 U3637 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b13), .B(n3395), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831792_127846048_127847952)
         );
  XOR2X1 U3638 ( .A(input_times_b0_mul_componentxUMxa2_and_b13), .B(n2459), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831792_127846048_127847952)
         );
  XOR2X1 U3639 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b12), .B(n2683), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831680_127845936_127847840)
         );
  XOR2X1 U3640 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b12), .B(n2917), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831680_127845936_127847840)
         );
  XOR2X1 U3641 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b12), .B(n3385), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831680_127845936_127847840)
         );
  XOR2X1 U3642 ( .A(input_times_b0_mul_componentxUMxa2_and_b12), .B(n2449), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831680_127845936_127847840)
         );
  XOR2X1 U3643 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b14), .B(n2703), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127831904_127846160_127848064)
         );
  XOR2X1 U3644 ( .A(input_times_b0_mul_componentxUMxa2_and_b14), .B(n2469), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127831904_127846160_127848064)
         );
  XOR2X1 U3645 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b7), .B(n2931), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127732816_127722496_127724400)
         );
  XOR2X1 U3646 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b7), .B(n3399), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127732816_127722496_127724400)
         );
  AND2X2 U3647 ( .A(input_p1_times_b1_mul_componentxUMxa1_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa0_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxcarry_layer1_127830168_127844480)
         );
  AND2X2 U3648 ( .A(input_p2_times_b2_mul_componentxUMxa1_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa0_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxcarry_layer1_127830168_127844480)
         );
  AND2X2 U3649 ( .A(output_p2_times_a2_mul_componentxUMxa1_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa0_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxcarry_layer1_127830168_127844480)
         );
  AND2X2 U3650 ( .A(input_times_b0_mul_componentxUMxa1_and_b0), 
        .B(input_times_b0_mul_componentxUMxa0_and_b1), 
        .Y(input_times_b0_mul_componentxUMxcarry_layer1_127830168_127844480)
         );
  XOR2X1 U3651 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127733040_127722720_127724624), 
        .B(n2777), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer2_128199368_128199480_128199648)
         );
  XOR2X1 U3652 ( 
        .A(input_p1_times_b1_mul_componentxUMxsum_layer1_127832016_127846272_127848176), 
        .B(input_p1_times_b1_mul_componentxUMxsum_layer1_127674016_127675920_127731136), 
        .Y(n2777) );
  XOR2X1 U3653 ( .A(input_p1_times_b1_mul_componentxUMxa8_and_b9), .B(n2715), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127733040_127722720_127724624)
         );
  XOR2X1 U3654 ( .A(input_p1_times_b1_mul_componentxUMxa2_and_b15), .B(n2713), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127832016_127846272_127848176)
         );
  XOR2X1 U3655 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127733040_127722720_127724624), 
        .B(n3011), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer2_128199368_128199480_128199648)
         );
  XOR2X1 U3656 ( 
        .A(input_p2_times_b2_mul_componentxUMxsum_layer1_127832016_127846272_127848176), 
        .B(input_p2_times_b2_mul_componentxUMxsum_layer1_127674016_127675920_127731136), 
        .Y(n3011) );
  XOR2X1 U3657 ( .A(input_p2_times_b2_mul_componentxUMxa8_and_b9), .B(n2949), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127733040_127722720_127724624)
         );
  XOR2X1 U3658 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b15), .B(n2947), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127832016_127846272_127848176)
         );
  XOR2X1 U3659 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127733040_127722720_127724624), 
        .B(n3479), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer2_128199368_128199480_128199648)
         );
  XOR2X1 U3660 ( 
        .A(output_p2_times_a2_mul_componentxUMxsum_layer1_127832016_127846272_127848176), 
        .B(output_p2_times_a2_mul_componentxUMxsum_layer1_127674016_127675920_127731136), 
        .Y(n3479) );
  XOR2X1 U3661 ( .A(output_p2_times_a2_mul_componentxUMxa8_and_b9), .B(n3417), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127733040_127722720_127724624)
         );
  XOR2X1 U3662 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b15), .B(n3415), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127832016_127846272_127848176)
         );
  XOR2X1 U3663 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127733040_127722720_127724624), 
        .B(n2543), 
        .Y(input_times_b0_mul_componentxUMxsum_layer2_128199368_128199480_128199648)
         );
  XOR2X1 U3664 ( 
        .A(input_times_b0_mul_componentxUMxsum_layer1_127832016_127846272_127848176), 
        .B(input_times_b0_mul_componentxUMxsum_layer1_127674016_127675920_127731136), 
        .Y(n2543) );
  XOR2X1 U3665 ( .A(input_times_b0_mul_componentxUMxa8_and_b9), .B(n2481), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127733040_127722720_127724624)
         );
  XOR2X1 U3666 ( .A(input_times_b0_mul_componentxUMxa2_and_b15), .B(n2479), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127832016_127846272_127848176)
         );
  INVX1 U3667 ( .A(n2930), .Y(n1038) );
  AOI22X1 U3668 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b11), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b12), .B0(n2929), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b10), .Y(n2930) );
  INVX1 U3669 ( .A(n3398), .Y(n561) );
  AOI22X1 U3670 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b11), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b12), .B0(n3397), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b10), .Y(n3398) );
  INVX1 U3671 ( .A(n2684), .Y(n919) );
  AOI22X1 U3672 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b13), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b14), .B0(n2683), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b12), .Y(n2684) );
  INVX1 U3673 ( .A(n2918), .Y(n1078) );
  AOI22X1 U3674 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b13), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b14), .B0(n2917), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b12), .Y(n2918) );
  INVX1 U3675 ( .A(n3386), .Y(n601) );
  AOI22X1 U3676 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b13), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b14), .B0(n3385), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b12), .Y(n3386) );
  INVX1 U3677 ( .A(n2450), .Y(n760) );
  AOI22X1 U3678 ( .A0(input_times_b0_mul_componentxUMxa1_and_b13), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b14), .B0(n2449), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b12), .Y(n2450) );
  INVX1 U3679 ( .A(n2694), .Y(n920) );
  AOI22X1 U3680 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b14), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b15), .B0(n2693), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b13), .Y(n2694) );
  INVX1 U3681 ( .A(n2928), .Y(n1079) );
  AOI22X1 U3682 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b14), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b15), .B0(n2927), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b13), .Y(n2928) );
  INVX1 U3683 ( .A(n3396), .Y(n602) );
  AOI22X1 U3684 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b14), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b15), .B0(n3395), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b13), .Y(n3396) );
  INVX1 U3685 ( .A(n2460), .Y(n761) );
  AOI22X1 U3686 ( .A0(input_times_b0_mul_componentxUMxa1_and_b14), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b15), .B0(n2459), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b13), .Y(n2460) );
  INVX1 U3687 ( .A(n2686), .Y(n887) );
  AOI22X1 U3688 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b10), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b11), .B0(n2685), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b9), .Y(n2686) );
  INVX1 U3689 ( .A(n2920), .Y(n1046) );
  AOI22X1 U3690 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b10), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b11), .B0(n2919), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b9), .Y(n2920) );
  INVX1 U3691 ( .A(n3388), .Y(n569) );
  AOI22X1 U3692 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b10), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b11), .B0(n3387), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b9), .Y(n3388) );
  INVX1 U3693 ( .A(n2452), .Y(n728) );
  AOI22X1 U3694 ( .A0(input_times_b0_mul_componentxUMxa4_and_b10), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b11), .B0(n2451), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b9), .Y(n2452) );
  INVX1 U3695 ( .A(n2698), .Y(n931) );
  AOI22X1 U3696 ( .A0(input_p1_times_b1_mul_componentxUMxa7_and_b8), 
        .A1(input_p1_times_b1_mul_componentxUMxa6_and_b9), .B0(n2697), 
        .B1(input_p1_times_b1_mul_componentxUMxa8_and_b7), .Y(n2698) );
  INVX1 U3697 ( .A(n2932), .Y(n1090) );
  AOI22X1 U3698 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b8), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b9), .B0(n2931), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b7), .Y(n2932) );
  INVX1 U3699 ( .A(n3400), .Y(n613) );
  AOI22X1 U3700 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b8), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b9), .B0(n3399), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b7), .Y(n3400) );
  INVX1 U3701 ( .A(n2464), .Y(n772) );
  AOI22X1 U3702 ( .A0(input_times_b0_mul_componentxUMxa7_and_b8), 
        .A1(input_times_b0_mul_componentxUMxa6_and_b9), .B0(n2463), 
        .B1(input_times_b0_mul_componentxUMxa8_and_b7), .Y(n2464) );
  INVX1 U3703 ( .A(n2706), .Y(n877) );
  AOI22X1 U3704 ( .A0(input_p1_times_b1_mul_componentxUMxa4_and_b12), 
        .A1(input_p1_times_b1_mul_componentxUMxa3_and_b13), .B0(n2705), 
        .B1(input_p1_times_b1_mul_componentxUMxa5_and_b11), .Y(n2706) );
  INVX1 U3705 ( .A(n2940), .Y(n1036) );
  AOI22X1 U3706 ( .A0(input_p2_times_b2_mul_componentxUMxa4_and_b12), 
        .A1(input_p2_times_b2_mul_componentxUMxa3_and_b13), .B0(n2939), 
        .B1(input_p2_times_b2_mul_componentxUMxa5_and_b11), .Y(n2940) );
  INVX1 U3707 ( .A(n3408), .Y(n559) );
  AOI22X1 U3708 ( .A0(output_p2_times_a2_mul_componentxUMxa4_and_b12), 
        .A1(output_p2_times_a2_mul_componentxUMxa3_and_b13), .B0(n3407), 
        .B1(output_p2_times_a2_mul_componentxUMxa5_and_b11), .Y(n3408) );
  INVX1 U3709 ( .A(n2472), .Y(n718) );
  AOI22X1 U3710 ( .A0(input_times_b0_mul_componentxUMxa4_and_b12), 
        .A1(input_times_b0_mul_componentxUMxa3_and_b13), .B0(n2471), 
        .B1(input_times_b0_mul_componentxUMxa5_and_b11), .Y(n2472) );
  INVX1 U3711 ( .A(n2942), .Y(n1081) );
  AOI22X1 U3712 ( .A0(input_p2_times_b2_mul_componentxUMxa7_and_b9), 
        .A1(input_p2_times_b2_mul_componentxUMxa6_and_b10), .B0(n2941), 
        .B1(input_p2_times_b2_mul_componentxUMxa8_and_b8), .Y(n2942) );
  INVX1 U3713 ( .A(n3410), .Y(n604) );
  AOI22X1 U3714 ( .A0(output_p2_times_a2_mul_componentxUMxa7_and_b9), 
        .A1(output_p2_times_a2_mul_componentxUMxa6_and_b10), .B0(n3409), 
        .B1(output_p2_times_a2_mul_componentxUMxa8_and_b8), .Y(n3410) );
  INVX1 U3715 ( .A(n2704), .Y(n921) );
  AOI22X1 U3716 ( .A0(input_p1_times_b1_mul_componentxUMxa1_and_b15), 
        .A1(input_p1_times_b1_mul_componentxUMxa0_and_b16), .B0(n2703), 
        .B1(input_p1_times_b1_mul_componentxUMxa2_and_b14), .Y(n2704) );
  INVX1 U3717 ( .A(n2938), .Y(n1080) );
  AOI22X1 U3718 ( .A0(input_p2_times_b2_mul_componentxUMxa1_and_b15), 
        .A1(input_p2_times_b2_mul_componentxUMxa0_and_b16), .B0(n2937), 
        .B1(input_p2_times_b2_mul_componentxUMxa2_and_b14), .Y(n2938) );
  INVX1 U3719 ( .A(n3406), .Y(n603) );
  AOI22X1 U3720 ( .A0(output_p2_times_a2_mul_componentxUMxa1_and_b15), 
        .A1(output_p2_times_a2_mul_componentxUMxa0_and_b16), .B0(n3405), 
        .B1(output_p2_times_a2_mul_componentxUMxa2_and_b14), .Y(n3406) );
  INVX1 U3721 ( .A(n2470), .Y(n762) );
  AOI22X1 U3722 ( .A0(input_times_b0_mul_componentxUMxa1_and_b15), 
        .A1(input_times_b0_mul_componentxUMxa0_and_b16), .B0(n2469), 
        .B1(input_times_b0_mul_componentxUMxa2_and_b14), .Y(n2470) );
  XOR2X1 U3723 ( .A(input_p1_times_b1_mul_componentxUMxa1_and_b0), 
        .B(input_p1_times_b1_mul_componentxUMxa0_and_b1), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[1]) );
  XOR2X1 U3724 ( .A(input_p2_times_b2_mul_componentxUMxa1_and_b0), 
        .B(input_p2_times_b2_mul_componentxUMxa0_and_b1), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[1]) );
  XOR2X1 U3725 ( .A(output_p2_times_a2_mul_componentxUMxa1_and_b0), 
        .B(output_p2_times_a2_mul_componentxUMxa0_and_b1), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[1]) );
  XOR2X1 U3726 ( .A(input_times_b0_mul_componentxUMxa1_and_b0), 
        .B(input_times_b0_mul_componentxUMxa0_and_b1), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[1]) );
  INVX1 U3727 ( .A(n4459), .Y(n995) );
  AOI22XL U3728 ( .A0(input_p1_times_b1_mul_componentxUMxfirst_vector[0]), 
        .A1(n125), .B0(input_p1_times_b1_mul_componentxUMxfirst_vector[0]), 
        .B1(n4442), .Y(n4459) );
  INVX1 U3729 ( .A(n4512), .Y(n1154) );
  AOI22XL U3730 ( .A0(input_p2_times_b2_mul_componentxUMxfirst_vector[0]), 
        .A1(n129), .B0(input_p2_times_b2_mul_componentxUMxfirst_vector[0]), 
        .B1(n4495), .Y(n4512) );
  INVX1 U3731 ( .A(n4618), .Y(n677) );
  AOI22XL U3732 ( .A0(output_p2_times_a2_mul_componentxUMxfirst_vector[0]), 
        .A1(n117), .B0(output_p2_times_a2_mul_componentxUMxfirst_vector[0]), 
        .B1(n4601), .Y(n4618) );
  INVX1 U3733 ( .A(input_times_b0_mul_componentxn108), .Y(n836) );
  AOI22XL U3734 ( .A0(input_times_b0_mul_componentxUMxfirst_vector[0]), 
        .A1(n121), .B0(input_times_b0_mul_componentxUMxfirst_vector[0]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn108) );
  XOR2X1 U3735 ( .A(n144), .B(n334), .Y(n81) );
  INVX1 U3736 ( .A(n81), .Y(n4442) );
  XOR2X1 U3737 ( .A(n142), .B(n325), .Y(n82) );
  INVX1 U3738 ( .A(n82), .Y(n4495) );
  XOR2X1 U3739 ( .A(n140), .B(n352), .Y(n83) );
  INVX1 U3740 ( .A(n83), .Y(n4601) );
  XOR2X1 U3741 ( .A(n132), .B(n343), .Y(n84) );
  INVX1 U3742 ( .A(n84), .Y(input_times_b0_mul_componentxn91) );
  XOR2X1 U3743 ( .A(input_p2_times_b2_mul_componentxUMxa2_and_b14), .B(n2937), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127831904_127846160_127848064)
         );
  XOR2X1 U3744 ( .A(output_p2_times_a2_mul_componentxUMxa2_and_b14), .B(n3405), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127831904_127846160_127848064)
         );
  INVX1 U3745 ( .A(n4450), .Y(n994) );
  AOI22X1 U3746 ( .A0(input_p1_times_b1_mul_componentxUMxfirst_vector[1]), 
        .A1(n126), 
        .B0(input_p1_times_b1_mul_componentxunsigned_output_inverted[1]), 
        .B1(n4442), .Y(n4450) );
  XOR2X1 U3747 ( .A(input_p1_times_b1_mul_componentxUMxfirst_vector[1]), 
        .B(input_p1_times_b1_mul_componentxUMxfirst_vector[0]), 
        .Y(input_p1_times_b1_mul_componentxunsigned_output_inverted[1]) );
  INVX1 U3748 ( .A(input_times_b0_mul_componentxn99), .Y(n835) );
  AOI22X1 U3749 ( .A0(input_times_b0_mul_componentxUMxfirst_vector[1]), 
        .A1(n122), 
        .B0(input_times_b0_mul_componentxunsigned_output_inverted[1]), 
        .B1(input_times_b0_mul_componentxn91), 
        .Y(input_times_b0_mul_componentxn99) );
  XOR2X1 U3750 ( .A(input_times_b0_mul_componentxUMxfirst_vector[1]), 
        .B(input_times_b0_mul_componentxUMxfirst_vector[0]), 
        .Y(input_times_b0_mul_componentxunsigned_output_inverted[1]) );
  INVX1 U3751 ( .A(n4503), .Y(n1153) );
  AOI22X1 U3752 ( .A0(input_p2_times_b2_mul_componentxUMxfirst_vector[1]), 
        .A1(n130), 
        .B0(input_p2_times_b2_mul_componentxunsigned_output_inverted[1]), 
        .B1(n4495), .Y(n4503) );
  XOR2X1 U3753 ( .A(input_p2_times_b2_mul_componentxUMxfirst_vector[1]), 
        .B(input_p2_times_b2_mul_componentxUMxfirst_vector[0]), 
        .Y(input_p2_times_b2_mul_componentxunsigned_output_inverted[1]) );
  INVX1 U3754 ( .A(n4609), .Y(n676) );
  AOI22X1 U3755 ( .A0(output_p2_times_a2_mul_componentxUMxfirst_vector[1]), 
        .A1(n118), 
        .B0(output_p2_times_a2_mul_componentxunsigned_output_inverted[1]), 
        .B1(n4601), .Y(n4609) );
  XOR2X1 U3756 ( .A(output_p2_times_a2_mul_componentxUMxfirst_vector[1]), 
        .B(output_p2_times_a2_mul_componentxUMxfirst_vector[0]), 
        .Y(output_p2_times_a2_mul_componentxunsigned_output_inverted[1]) );
  OAI2BB2X1 U3757 ( .B0(n131), .B1(n319), .A0N(input_previous_1[17]), 
        .A1N(n321), .Y(n4636) );
  OAI2BB2X1 U3758 ( .B0(n143), .B1(n319), .A0N(input_previous_2[17]), 
        .A1N(n320), .Y(n4654) );
  NAND3BX1 U3759 ( .AN(n845), .B(input_times_b0_div_componentxn54), 
        .C(input_times_b0_div_componentxUDxinverter_for_substractionxn2), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn16) );
  NAND3BX1 U3760 ( .AN(n1004), .B(n4232), .C(n1761), .Y(n1768) );
  NAND3BX1 U3761 ( .AN(n1163), .B(n4288), .C(n1770), .Y(n1777) );
  NAND3BX1 U3762 ( .AN(n527), .B(n4342), .C(n1779), .Y(n1786) );
  NAND3BX1 U3763 ( .AN(n686), .B(n4398), .C(n1788), .Y(n1795) );
  NOR2BX1 U3764 ( .AN(n3892), .B(\parameter_B0_div[7] ), .Y(n3891) );
  NOR2BX1 U3765 ( .AN(n3935), .B(\parameter_B1_div[7] ), .Y(n3934) );
  NOR2BX1 U3766 ( .AN(n3978), .B(\parameter_B2_div[7] ), .Y(n3977) );
  NOR2BX1 U3767 ( .AN(n4021), .B(\parameter_A1_div[7] ), .Y(n4020) );
  NOR2BX1 U3768 ( .AN(n4064), .B(\parameter_A2_div[7] ), .Y(n4063) );
  NOR2X1 U3769 ( .A(\parameter_B0_div[7] ), .B(n3893), .Y(n3892) );
  NOR2X1 U3770 ( .A(\parameter_B1_div[7] ), .B(n3936), .Y(n3935) );
  NOR2X1 U3771 ( .A(\parameter_B2_div[7] ), .B(n3979), .Y(n3978) );
  NOR2X1 U3772 ( .A(\parameter_A1_div[7] ), .B(n4022), .Y(n4021) );
  NOR2X1 U3773 ( .A(\parameter_A2_div[7] ), .B(n4065), .Y(n4064) );
  XOR2X1 U3774 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn2), 
        .B(input_times_b0_div_componentxn54), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[9]) );
  XOR2X1 U3775 ( .A(n1761), .B(n4232), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[9])
         );
  XOR2X1 U3776 ( .A(n1770), .B(n4288), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[9])
         );
  XOR2X1 U3777 ( .A(n1779), .B(n4342), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[9])
         );
  XOR2X1 U3778 ( .A(n1788), .B(n4398), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[9])
         );
  XOR2X1 U3779 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn8), 
        .B(n849), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[3]) );
  XOR2X1 U3780 ( .A(n1764), .B(n1008), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[3])
         );
  XOR2X1 U3781 ( .A(n1773), .B(n1167), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[3])
         );
  XOR2X1 U3782 ( .A(n1782), .B(n531), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[3])
         );
  XOR2X1 U3783 ( .A(n1791), .B(n690), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[3])
         );
  XOR2X1 U3784 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn6), 
        .B(n851), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[5]) );
  XOR2X1 U3785 ( .A(n1763), .B(n1010), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[5])
         );
  XOR2X1 U3786 ( .A(n1772), .B(n1169), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[5])
         );
  XOR2X1 U3787 ( .A(n1781), .B(n533), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[5])
         );
  XOR2X1 U3788 ( .A(n1790), .B(n692), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[5])
         );
  OR3XL U3789 ( .A(n851), .B(n852), 
        .C(input_times_b0_div_componentxUDxinverter_for_substractionxn6), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn4) );
  OR3XL U3790 ( .A(n1010), .B(n1011), .C(n1763), .Y(n1762) );
  OR3XL U3791 ( .A(n1169), .B(n1170), .C(n1772), .Y(n1771) );
  OR3XL U3792 ( .A(n533), .B(n534), .C(n1781), .Y(n1780) );
  OR3XL U3793 ( .A(n692), .B(n693), .C(n1790), .Y(n1789) );
  OR2X2 U3794 ( .A(n3895), .B(\parameter_B0_div[7] ), .Y(n3893) );
  OR2X2 U3795 ( .A(n3938), .B(\parameter_B1_div[7] ), .Y(n3936) );
  OR2X2 U3796 ( .A(n3981), .B(\parameter_B2_div[7] ), .Y(n3979) );
  OR2X2 U3797 ( .A(n4024), .B(\parameter_A1_div[7] ), .Y(n4022) );
  OR2X2 U3798 ( .A(n4067), .B(\parameter_A2_div[7] ), .Y(n4065) );
  XNOR2X1 U3799 ( .A(n85), .B(n850), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[4]) );
  NOR2X1 U3800 ( .A(n849), 
        .B(input_times_b0_div_componentxUDxinverter_for_substractionxn8), 
        .Y(n85) );
  XNOR2X1 U3801 ( .A(n86), .B(n1009), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[4])
         );
  NOR2X1 U3802 ( .A(n1008), .B(n1764), .Y(n86) );
  XNOR2X1 U3803 ( .A(n87), .B(n1168), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[4])
         );
  NOR2X1 U3804 ( .A(n1167), .B(n1773), .Y(n87) );
  XNOR2X1 U3805 ( .A(n88), .B(n532), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[4])
         );
  NOR2X1 U3806 ( .A(n531), .B(n1782), .Y(n88) );
  XNOR2X1 U3807 ( .A(n89), .B(n691), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[4])
         );
  NOR2X1 U3808 ( .A(n690), .B(n1791), .Y(n89) );
  XNOR2X1 U3809 ( .A(n90), .B(n852), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[6]) );
  NOR2X1 U3810 ( .A(n851), 
        .B(input_times_b0_div_componentxUDxinverter_for_substractionxn6), 
        .Y(n90) );
  XNOR2X1 U3811 ( .A(n91), .B(n1011), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[6])
         );
  NOR2X1 U3812 ( .A(n1010), .B(n1763), .Y(n91) );
  XNOR2X1 U3813 ( .A(n92), .B(n1170), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[6])
         );
  NOR2X1 U3814 ( .A(n1169), .B(n1772), .Y(n92) );
  XNOR2X1 U3815 ( .A(n93), .B(n534), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[6])
         );
  NOR2X1 U3816 ( .A(n533), .B(n1781), .Y(n93) );
  XNOR2X1 U3817 ( .A(n94), .B(n693), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[6])
         );
  NOR2X1 U3818 ( .A(n692), .B(n1790), .Y(n94) );
  XOR2X1 U3819 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn18), 
        .B(n845), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[10]) );
  NAND2X1 U3820 ( 
        .A(input_times_b0_div_componentxUDxinverter_for_substractionxn2), 
        .B(input_times_b0_div_componentxn54), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn18) );
  XOR2X1 U3821 ( .A(n1769), .B(n1004), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[10])
         );
  NAND2X1 U3822 ( .A(n1761), .B(n4232), .Y(n1769) );
  XOR2X1 U3823 ( .A(n1778), .B(n1163), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[10])
         );
  NAND2X1 U3824 ( .A(n1770), .B(n4288), .Y(n1778) );
  XOR2X1 U3825 ( .A(n1787), .B(n527), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[10])
         );
  NAND2X1 U3826 ( .A(n1779), .B(n4342), .Y(n1787) );
  XOR2X1 U3827 ( .A(n1796), .B(n686), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[10])
         );
  NAND2X1 U3828 ( .A(n1788), .B(n4398), .Y(n1796) );
  OR3XL U3829 ( .A(n849), .B(n850), 
        .C(input_times_b0_div_componentxUDxinverter_for_substractionxn8), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn6) );
  OR3XL U3830 ( .A(n1008), .B(n1009), .C(n1764), .Y(n1763) );
  OR3XL U3831 ( .A(n1167), .B(n1168), .C(n1773), .Y(n1772) );
  OR3XL U3832 ( .A(n531), .B(n532), .C(n1782), .Y(n1781) );
  OR3XL U3833 ( .A(n690), .B(n691), .C(n1791), .Y(n1790) );
  INVX1 U3834 ( .A(input_times_b0_div_componentxn52), .Y(n853) );
  INVX1 U3835 ( .A(n4230), .Y(n1012) );
  INVX1 U3836 ( .A(n4286), .Y(n1171) );
  INVX1 U3837 ( .A(n4340), .Y(n535) );
  INVX1 U3838 ( .A(n4396), .Y(n694) );
  INVX1 U3839 ( .A(input_times_b0_div_componentxn58), .Y(n840) );
  INVX1 U3840 ( .A(n4236), .Y(n999) );
  INVX1 U3841 ( .A(n4292), .Y(n1158) );
  INVX1 U3842 ( .A(n4346), .Y(n522) );
  INVX1 U3843 ( .A(n4402), .Y(n681) );
  INVX1 U3844 ( .A(input_times_b0_div_componentxn56), .Y(n838) );
  INVX1 U3845 ( .A(n4234), .Y(n997) );
  INVX1 U3846 ( .A(n4290), .Y(n1156) );
  INVX1 U3847 ( .A(n4344), .Y(n520) );
  INVX1 U3848 ( .A(n4400), .Y(n679) );
  INVX1 U3849 ( .A(input_times_b0_div_componentxn53), .Y(n854) );
  INVX1 U3850 ( .A(n4231), .Y(n1013) );
  INVX1 U3851 ( .A(n4287), .Y(n1172) );
  INVX1 U3852 ( .A(n4341), .Y(n536) );
  INVX1 U3853 ( .A(n4397), .Y(n695) );
  XNOR2X1 U3854 ( .A(n95), .B(n843), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[16]) );
  NOR2X1 U3855 ( .A(n842), 
        .B(input_times_b0_div_componentxUDxinverter_for_substractionxn12), 
        .Y(n95) );
  XNOR2X1 U3856 ( .A(n96), .B(n1002), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[16])
         );
  NOR2X1 U3857 ( .A(n1001), .B(n1766), .Y(n96) );
  XNOR2X1 U3858 ( .A(n97), .B(n1161), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[16])
         );
  NOR2X1 U3859 ( .A(n1160), .B(n1775), .Y(n97) );
  XNOR2X1 U3860 ( .A(n98), .B(n525), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[16])
         );
  NOR2X1 U3861 ( .A(n524), .B(n1784), .Y(n98) );
  XNOR2X1 U3862 ( .A(n99), .B(n684), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[16])
         );
  NOR2X1 U3863 ( .A(n683), .B(n1793), .Y(n99) );
  INVX1 U3864 ( .A(input_times_b0_div_componentxn57), .Y(n839) );
  INVX1 U3865 ( .A(n4235), .Y(n998) );
  INVX1 U3866 ( .A(n4291), .Y(n1157) );
  INVX1 U3867 ( .A(n4345), .Y(n521) );
  INVX1 U3868 ( .A(n4401), .Y(n680) );
  INVX1 U3869 ( .A(input_times_b0_div_componentxn59), .Y(n841) );
  INVX1 U3870 ( .A(n4237), .Y(n1000) );
  INVX1 U3871 ( .A(n4293), .Y(n1159) );
  INVX1 U3872 ( .A(n4347), .Y(n523) );
  INVX1 U3873 ( .A(n4403), .Y(n682) );
  INVX1 U3874 ( .A(input_times_b0_div_componentxn55), .Y(n845) );
  INVX1 U3875 ( .A(n4233), .Y(n1004) );
  INVX1 U3876 ( .A(n4289), .Y(n1163) );
  INVX1 U3877 ( .A(n4343), .Y(n527) );
  INVX1 U3878 ( .A(n4399), .Y(n686) );
  INVX1 U3879 ( .A(input_times_b0_div_componentxn60), .Y(n842) );
  INVX1 U3880 ( .A(n4238), .Y(n1001) );
  INVX1 U3881 ( .A(n4294), .Y(n1160) );
  INVX1 U3882 ( .A(n4348), .Y(n524) );
  INVX1 U3883 ( .A(n4404), .Y(n683) );
  INVX1 U3884 ( .A(n317), .Y(n291) );
  INVX1 U3885 ( .A(n317), .Y(n292) );
  INVX1 U3886 ( .A(n317), .Y(n293) );
  INVX1 U3887 ( .A(n316), .Y(n294) );
  INVX1 U3888 ( .A(n316), .Y(n295) );
  INVX1 U3889 ( .A(n316), .Y(n296) );
  INVX1 U3890 ( .A(n317), .Y(n297) );
  INVX1 U3891 ( .A(reset), .Y(n284) );
  INVX1 U3892 ( .A(n318), .Y(n285) );
  INVX1 U3893 ( .A(n315), .Y(n286) );
  INVX1 U3894 ( .A(n315), .Y(n287) );
  INVX1 U3895 ( .A(n318), .Y(n288) );
  INVX1 U3896 ( .A(n318), .Y(n289) );
  INVX1 U3897 ( .A(n318), .Y(n290) );
  INVX1 U3898 ( .A(reset), .Y(n307) );
  INVX1 U3899 ( .A(reset), .Y(n308) );
  INVX1 U3900 ( .A(n317), .Y(n309) );
  INVX1 U3901 ( .A(n316), .Y(n310) );
  INVX1 U3902 ( .A(n318), .Y(n311) );
  INVX1 U3903 ( .A(n315), .Y(n312) );
  INVX1 U3904 ( .A(n315), .Y(n313) );
  INVX1 U3905 ( .A(n316), .Y(n298) );
  INVX1 U3906 ( .A(n318), .Y(n299) );
  INVX1 U3907 ( .A(n318), .Y(n300) );
  INVX1 U3908 ( .A(reset), .Y(n301) );
  INVX1 U3909 ( .A(n315), .Y(n302) );
  INVX1 U3910 ( .A(n317), .Y(n303) );
  INVX1 U3911 ( .A(n316), .Y(n304) );
  INVX1 U3912 ( .A(n316), .Y(n305) );
  INVX1 U3913 ( .A(n317), .Y(n306) );
  INVX1 U3914 ( .A(reset), .Y(n283) );
  INVX1 U3915 ( .A(n315), .Y(n314) );
  AOI32X1 U3916 ( .A0(n1320), .A1(n4135), .A2(n1340), .B0(n1311), .B1(n1331), 
        .Y(n4134) );
  AOI32X1 U3917 ( .A0(n1379), .A1(results_b0_b1_adderxn19), .A2(n1237), 
        .B0(n1370), .B1(n1227), .Y(results_b0_b1_adderxn17) );
  AOI22X1 U3918 ( .A0(n1309), .A1(n1329), .B0(n4131), .B1(n4132), .Y(n4130) );
  AOI22X1 U3919 ( .A0(n1368), .A1(n1223), .B0(results_b0_b1_adderxn14), 
        .B1(results_b0_b1_adderxn15), .Y(results_b0_b1_adderxn13) );
  AOI22X1 U3920 ( .A0(n1307), .A1(n1327), .B0(n4127), .B1(n4128), .Y(n4126) );
  AOI22X1 U3921 ( .A0(n1348), .A1(results_b0_b1[3]), .B0(n4098), .B1(n4099), 
        .Y(n4097) );
  AOI22X1 U3922 ( .A0(n1366), .A1(n1219), .B0(results_b0_b1_adderxn10), 
        .B1(results_b0_b1_adderxn11), .Y(results_b0_b1_adderxn9) );
  AOI22X1 U3923 ( .A0(n1305), .A1(n1325), .B0(n4123), .B1(n4124), .Y(n4122) );
  AOI22X1 U3924 ( .A0(n1346), .A1(results_b0_b1[5]), .B0(n4094), .B1(n4095), 
        .Y(n4093) );
  AOI22X1 U3925 ( .A0(n1364), .A1(n1215), .B0(results_b0_b1_adderxn6), 
        .B1(results_b0_b1_adderxn7), .Y(results_b0_b1_adderxn5) );
  AOI22X1 U3926 ( .A0(n1344), .A1(results_b0_b1[7]), .B0(n4090), .B1(n4091), 
        .Y(n4089) );
  AOI22X1 U3927 ( .A0(n1362), .A1(n1211), .B0(results_b0_b1_adderxn2), 
        .B1(results_b0_b1_adderxn3), .Y(results_b0_b1_adderxn34) );
  AOI22X1 U3928 ( .A0(n1342), .A1(results_b0_b1[9]), .B0(n4086), .B1(n4087), 
        .Y(n4117) );
  AOI22X1 U3929 ( .A0(n1377), .A1(n1234), .B0(results_b0_b1_adderxn32), 
        .B1(results_b0_b1_adderxn33), .Y(results_b0_b1_adderxn30) );
  AOI22X1 U3930 ( .A0(n1357), .A1(results_b0_b1[11]), .B0(n4115), .B1(n4116), 
        .Y(n4113) );
  AOI22X1 U3931 ( .A0(n1375), .A1(n1232), .B0(results_b0_b1_adderxn28), 
        .B1(results_b0_b1_adderxn29), .Y(results_b0_b1_adderxn26) );
  AOI22X1 U3932 ( .A0(n1355), .A1(results_b0_b1[13]), .B0(n4111), .B1(n4112), 
        .Y(n4109) );
  OAI2BB2X1 U3933 ( .B0(n4101), .B1(n4100), .A0N(n1349), 
        .A1N(results_b0_b1[2]), .Y(n4098) );
  OAI2BB2X1 U3934 ( .B0(n4134), .B1(n4133), .A0N(n1310), .A1N(n1330), 
        .Y(n4131) );
  OAI2BB2X1 U3935 ( .B0(results_b0_b1_adderxn17), .B1(results_b0_b1_adderxn16), 
        .A0N(n1369), .A1N(n1225), .Y(results_b0_b1_adderxn14) );
  OAI2BB2X1 U3936 ( .B0(n4130), .B1(n4129), .A0N(n1308), .A1N(n1328), 
        .Y(n4127) );
  OAI2BB2X1 U3937 ( .B0(results_b0_b1_adderxn13), .B1(results_b0_b1_adderxn12), 
        .A0N(n1367), .A1N(n1221), .Y(results_b0_b1_adderxn10) );
  OAI2BB2X1 U3938 ( .B0(n4097), .B1(n4096), .A0N(n1347), 
        .A1N(results_b0_b1[4]), .Y(n4094) );
  OAI2BB2X1 U3939 ( .B0(n4126), .B1(n4125), .A0N(n1306), .A1N(n1326), 
        .Y(n4123) );
  OAI2BB2X1 U3940 ( .B0(results_b0_b1_adderxn9), .B1(results_b0_b1_adderxn8), 
        .A0N(n1365), .A1N(n1217), .Y(results_b0_b1_adderxn6) );
  OAI2BB2X1 U3941 ( .B0(n4093), .B1(n4092), .A0N(n1345), 
        .A1N(results_b0_b1[6]), .Y(n4090) );
  OAI2BB2X1 U3942 ( .B0(results_b0_b1_adderxn5), .B1(results_b0_b1_adderxn4), 
        .A0N(n1363), .A1N(n1213), .Y(results_b0_b1_adderxn2) );
  OAI2BB2X1 U3943 ( .B0(n4089), .B1(n4088), .A0N(n1343), 
        .A1N(results_b0_b1[8]), .Y(n4086) );
  OAI2BB2X1 U3944 ( .B0(results_b0_b1_adderxn34), .B1(results_b0_b1_adderxn35), 
        .A0N(n1378), .A1N(n1235), .Y(results_b0_b1_adderxn32) );
  OAI2BB2X1 U3945 ( .B0(n4117), .B1(n4118), .A0N(n1358), 
        .A1N(results_b0_b1[10]), .Y(n4115) );
  OAI2BB2X1 U3946 ( .B0(results_b0_b1_adderxn30), .B1(results_b0_b1_adderxn31), 
        .A0N(n1376), .A1N(n1233), .Y(results_b0_b1_adderxn28) );
  OAI2BB2X1 U3947 ( .B0(n4113), .B1(n4114), .A0N(n1356), 
        .A1N(results_b0_b1[12]), .Y(n4111) );
  OAI2BB2X1 U3948 ( .B0(n4109), .B1(n4110), .A0N(n1354), 
        .A1N(results_b0_b1[14]), .Y(n4107) );
  NOR2X1 U3949 ( .A(n218), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b3) );
  NOR2X1 U3950 ( .A(n217), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b4) );
  NOR2X1 U3951 ( .A(n231), .B(n216), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b5) );
  XOR2X1 U3952 ( .A(results_b0_b1[3]), .B(n1348), .Y(n4099) );
  XOR2X1 U3953 ( .A(results_b0_b1[5]), .B(n1346), .Y(n4095) );
  XOR2X1 U3954 ( .A(results_b0_b1[7]), .B(n1344), .Y(n4091) );
  XOR2X1 U3955 ( .A(results_b0_b1[9]), .B(n1342), .Y(n4087) );
  XOR2X1 U3956 ( .A(results_b0_b1[11]), .B(n1357), .Y(n4116) );
  XOR2X1 U3957 ( .A(results_b0_b1[13]), .B(n1355), .Y(n4112) );
  XOR2X1 U3958 ( .A(n1331), .B(n1311), .Y(n4135) );
  XOR2X1 U3959 ( .A(n1227), .B(n1370), .Y(results_b0_b1_adderxn19) );
  XNOR2X1 U3960 ( .A(results_b0_b1[2]), .B(n1349), .Y(n4100) );
  XNOR2X1 U3961 ( .A(results_b0_b1[4]), .B(n1347), .Y(n4096) );
  XNOR2X1 U3962 ( .A(results_b0_b1[6]), .B(n1345), .Y(n4092) );
  XNOR2X1 U3963 ( .A(results_b0_b1[8]), .B(n1343), .Y(n4088) );
  XNOR2X1 U3964 ( .A(results_b0_b1[10]), .B(n1358), .Y(n4118) );
  XNOR2X1 U3965 ( .A(results_b0_b1[12]), .B(n1356), .Y(n4114) );
  XNOR2X1 U3966 ( .A(results_b0_b1[14]), .B(n1354), .Y(n4110) );
  INVX1 U3967 ( .A(n169), .Y(n1321) );
  INVX1 U3968 ( .A(n168), .Y(n1341) );
  INVX1 U3969 ( .A(n166), .Y(n1380) );
  INVX1 U3970 ( .A(n260), .Y(n1238) );
  AOI32X1 U3971 ( .A0(n1359), .A1(n4102), .A2(results_b0_b1[0]), .B0(n1350), 
        .B1(results_b0_b1[1]), .Y(n4101) );
  AOI22X1 U3972 ( .A0(n1303), .A1(n1323), .B0(n4119), .B1(n4120), .Y(n4150) );
  AOI22X1 U3973 ( .A0(n1318), .A1(n1338), .B0(n4148), .B1(n4149), .Y(n4146) );
  AOI22X1 U3974 ( .A0(n1316), .A1(n1336), .B0(n4144), .B1(n4145), .Y(n4142) );
  XOR2X1 U3975 ( .A(n1320), .B(n1340), .Y(results_a1_a2_inv[0]) );
  NOR2X1 U3976 ( .A(n220), .B(n4545), 
        .Y(output_p1_times_a1_mul_componentxUMxa10_and_b1) );
  NOR2X1 U3977 ( .A(n219), .B(n4545), 
        .Y(output_p1_times_a1_mul_componentxUMxa10_and_b2) );
  OAI2BB2X1 U3978 ( .B0(n4122), .B1(n4121), .A0N(n1304), .A1N(n1324), 
        .Y(n4119) );
  OAI2BB2X1 U3979 ( .B0(n4150), .B1(n4151), .A0N(n1319), .A1N(n1339), 
        .Y(n4148) );
  OAI2BB2X1 U3980 ( .B0(n4146), .B1(n4147), .A0N(n1317), .A1N(n1337), 
        .Y(n4144) );
  OAI2BB2X1 U3981 ( .B0(results_b0_b1_adderxn26), .B1(results_b0_b1_adderxn27), 
        .A0N(n1374), .A1N(n1231), .Y(results_b0_b1_adderxn24) );
  OAI2BB2X1 U3982 ( .B0(n4142), .B1(n4143), .A0N(n1315), .A1N(n1335), 
        .Y(n4140) );
  NOR2X1 U3983 ( .A(n220), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b1) );
  NOR2X1 U3984 ( .A(n220), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b1) );
  NOR2X1 U3985 ( .A(n220), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b1) );
  NOR2X1 U3986 ( .A(n219), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b2) );
  NOR2X1 U3987 ( .A(n219), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b2) );
  NOR2X1 U3988 ( .A(n219), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b2) );
  NOR2X1 U3989 ( .A(n218), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b3) );
  NOR2X1 U3990 ( .A(n218), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b3) );
  NOR2X1 U3991 ( .A(n217), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b4) );
  NOR2X1 U3992 ( .A(n217), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b4) );
  NOR2X1 U3993 ( .A(n216), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b5) );
  NOR2X1 U3994 ( .A(n216), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b5) );
  NOR2X1 U3995 ( .A(n216), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b5) );
  NOR2X1 U3996 ( .A(n215), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b6) );
  NOR2X1 U3997 ( .A(n215), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b6) );
  AOI22X1 U3998 ( .A0(n4138), .A1(n1301), .B0(n1333), .B1(n1313), .Y(n4137) );
  NOR2X1 U3999 ( .A(n221), .B(n4544), 
        .Y(output_p1_times_a1_mul_componentxUMxa11_and_b0) );
  NOR2X1 U4000 ( .A(n231), .B(n217), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b4) );
  NOR2X1 U4001 ( .A(n231), .B(n218), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b3) );
  NOR2X1 U4002 ( .A(n231), .B(n219), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b2) );
  NOR2X1 U4003 ( .A(n231), .B(n215), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b6) );
  NOR2X1 U4004 ( .A(n221), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b0) );
  NOR2X1 U4005 ( .A(n219), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b2) );
  NOR2X1 U4006 ( .A(n219), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b2) );
  NOR2X1 U4007 ( .A(n218), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b3) );
  NOR2X1 U4008 ( .A(n218), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b3) );
  NOR2X1 U4009 ( .A(n217), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b4) );
  NOR2X1 U4010 ( .A(n217), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b4) );
  NOR2X1 U4011 ( .A(n216), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b5) );
  NOR2X1 U4012 ( .A(n216), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b5) );
  NOR2X1 U4013 ( .A(n215), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b6) );
  NOR2X1 U4014 ( .A(n215), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b6) );
  NOR2X1 U4015 ( .A(n222), .B(n219), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b2) );
  NOR2X1 U4016 ( .A(n221), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b0) );
  NOR2X1 U4017 ( .A(n221), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b0) );
  NOR2X1 U4018 ( .A(n220), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b1) );
  NOR2X1 U4019 ( .A(n220), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b1) );
  NOR2X1 U4020 ( .A(n219), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b2) );
  NOR2X1 U4021 ( .A(n219), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b2) );
  NOR2X1 U4022 ( .A(n218), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b3) );
  NOR2X1 U4023 ( .A(n218), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b3) );
  NOR2X1 U4024 ( .A(n217), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b4) );
  NOR2X1 U4025 ( .A(n217), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b4) );
  NOR2X1 U4026 ( .A(n216), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b5) );
  NOR2X1 U4027 ( .A(n216), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b5) );
  NOR2X1 U4028 ( .A(n215), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b6) );
  NOR2X1 U4029 ( .A(n220), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b1) );
  NOR2X1 U4030 ( .A(n220), .B(n225), 
        .Y(output_p1_times_a1_mul_componentxUMxa6_and_b1) );
  NOR2X1 U4031 ( .A(n221), .B(n227), 
        .Y(output_p1_times_a1_mul_componentxUMxa4_and_b0) );
  NOR2X1 U4032 ( .A(n221), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b0) );
  XOR2X1 U4033 ( .A(n1359), .B(results_b0_b1[0]), .Y(results_b0_b1_b2[0]) );
  XOR2X1 U4034 ( .A(n1379), .B(n1237), .Y(results_b0_b1[0]) );
  XOR2X1 U4035 ( .A(n1329), .B(n1309), .Y(n4132) );
  XOR2X1 U4036 ( .A(n1223), .B(n1368), .Y(results_b0_b1_adderxn15) );
  XOR2X1 U4037 ( .A(n1327), .B(n1307), .Y(n4128) );
  XOR2X1 U4038 ( .A(n1219), .B(n1366), .Y(results_b0_b1_adderxn11) );
  XOR2X1 U4039 ( .A(n1325), .B(n1305), .Y(n4124) );
  XOR2X1 U4040 ( .A(n1215), .B(n1364), .Y(results_b0_b1_adderxn7) );
  XOR2X1 U4041 ( .A(n1323), .B(n1303), .Y(n4120) );
  XOR2X1 U4042 ( .A(n1211), .B(n1362), .Y(results_b0_b1_adderxn3) );
  XOR2X1 U4043 ( .A(n1234), .B(n1377), .Y(results_b0_b1_adderxn33) );
  XOR2X1 U4044 ( .A(n1232), .B(n1375), .Y(results_b0_b1_adderxn29) );
  XOR2X1 U4045 ( .A(results_b0_b1[15]), .B(n1353), .Y(n4108) );
  XNOR2X1 U4046 ( .A(n100), .B(n4135), .Y(results_a1_a2[1]) );
  NAND2X1 U4047 ( .A(n1340), .B(n1320), .Y(n100) );
  XOR2X1 U4048 ( .A(results_b0_b1[1]), .B(n1350), .Y(n4102) );
  XNOR2X1 U4049 ( .A(n1330), .B(n1310), .Y(n4133) );
  XNOR2X1 U4050 ( .A(n1225), .B(n1369), .Y(results_b0_b1_adderxn16) );
  XNOR2X1 U4051 ( .A(n1328), .B(n1308), .Y(n4129) );
  XNOR2X1 U4052 ( .A(n1221), .B(n1367), .Y(results_b0_b1_adderxn12) );
  XNOR2X1 U4053 ( .A(n1326), .B(n1306), .Y(n4125) );
  XNOR2X1 U4054 ( .A(n1217), .B(n1365), .Y(results_b0_b1_adderxn8) );
  XNOR2X1 U4055 ( .A(n1324), .B(n1304), .Y(n4121) );
  XNOR2X1 U4056 ( .A(n1213), .B(n1363), .Y(results_b0_b1_adderxn4) );
  XNOR2X1 U4057 ( .A(n1235), .B(n1378), .Y(results_b0_b1_adderxn35) );
  XNOR2X1 U4058 ( .A(n1233), .B(n1376), .Y(results_b0_b1_adderxn31) );
  XNOR2X1 U4059 ( .A(n1231), .B(n1374), .Y(results_b0_b1_adderxn27) );
  XOR2X1 U4060 ( .A(results_b0_b1[16]), .B(n1352), .Y(n4105) );
  XNOR2X1 U4061 ( .A(n101), .B(results_b0_b1_adderxn19), .Y(results_b0_b1[1])
         );
  NAND2X1 U4062 ( .A(n1237), .B(n1379), .Y(n101) );
  XNOR2X1 U4063 ( .A(n102), .B(n4102), .Y(results_b0_b1_b2[1]) );
  NAND2X1 U4064 ( .A(results_b0_b1[0]), .B(n1359), .Y(n102) );
  XOR2X1 U4065 ( .A(results_a1_a2_inv_inverterxn10), .B(results_a1_a2[17]), 
        .Y(results_a1_a2_inv[17]) );
  NAND2BX1 U4066 ( .AN(results_a1_a2[16]), .B(results_a1_a2_inv_inverterxn11), 
        .Y(results_a1_a2_inv_inverterxn10) );
  XOR2X1 U4067 ( .A(n4136), .B(n4137), .Y(results_a1_a2[17]) );
  XNOR2X1 U4068 ( .A(n1312), .B(n1332), .Y(n4136) );
  XOR2X1 U4069 ( .A(results_b0_b1_adderxn20), .B(results_b0_b1_adderxn21), 
        .Y(results_b0_b1[17]) );
  XNOR2X1 U4070 ( .A(n1371), .B(n1228), .Y(results_b0_b1_adderxn20) );
  AOI22X1 U4071 ( .A0(results_b0_b1_adderxn22), .A1(n1209), .B0(n1229), 
        .B1(n1372), .Y(results_b0_b1_adderxn21) );
  INVX1 U4072 ( .A(n4194), .Y(n1371) );
  XOR2X1 U4073 ( .A(n4103), .B(n4104), .Y(results_b0_b1_b2[17]) );
  XNOR2X1 U4074 ( .A(n1351), .B(results_b0_b1[17]), .Y(n4103) );
  AOI22X1 U4075 ( .A0(n4105), .A1(n1207), .B0(results_b0_b1[16]), .B1(n1352), 
        .Y(n4104) );
  INVX1 U4076 ( .A(n4250), .Y(n1351) );
  INVX1 U4077 ( .A(n167), .Y(n1360) );
  XNOR2X1 U4078 ( .A(n112), .B(n360), .Y(n4315) );
  INVX1 U4079 ( .A(results_b0_b1_adderxn23), .Y(n1209) );
  AOI22X1 U4080 ( .A0(n1373), .A1(n1230), .B0(results_b0_b1_adderxn24), 
        .B1(results_b0_b1_adderxn25), .Y(results_b0_b1_adderxn23) );
  INVX1 U4081 ( .A(n4139), .Y(n1301) );
  AOI22X1 U4082 ( .A0(n1314), .A1(n1334), .B0(n4140), .B1(n4141), .Y(n4139) );
  INVX1 U4083 ( .A(n4106), .Y(n1207) );
  AOI22X1 U4084 ( .A0(n1353), .A1(results_b0_b1[15]), .B0(n4107), .B1(n4108), 
        .Y(n4106) );
  NOR2X1 U4085 ( .A(n218), .B(n4545), 
        .Y(output_p1_times_a1_mul_componentxUMxa10_and_b3) );
  NOR2X1 U4086 ( .A(n217), .B(n4545), 
        .Y(output_p1_times_a1_mul_componentxUMxa10_and_b4) );
  NOR2X1 U4087 ( .A(n220), .B(n4542), 
        .Y(output_p1_times_a1_mul_componentxUMxa13_and_b1) );
  NOR2X1 U4088 ( .A(n219), .B(n4542), 
        .Y(output_p1_times_a1_mul_componentxUMxa13_and_b2) );
  NOR2X1 U4089 ( .A(n215), .B(n224), 
        .Y(output_p1_times_a1_mul_componentxUMxa7_and_b6) );
  NOR2X1 U4090 ( .A(n220), .B(n4544), 
        .Y(output_p1_times_a1_mul_componentxUMxa11_and_b1) );
  NOR2X1 U4091 ( .A(n219), .B(n4544), 
        .Y(output_p1_times_a1_mul_componentxUMxa11_and_b2) );
  NOR2X1 U4092 ( .A(n218), .B(n4544), 
        .Y(output_p1_times_a1_mul_componentxUMxa11_and_b3) );
  NOR2X1 U4093 ( .A(n221), .B(n4543), 
        .Y(output_p1_times_a1_mul_componentxUMxa12_and_b0) );
  NOR2X1 U4094 ( .A(n219), .B(n4543), 
        .Y(output_p1_times_a1_mul_componentxUMxa12_and_b2) );
  NOR2X1 U4095 ( .A(n220), .B(n4543), 
        .Y(output_p1_times_a1_mul_componentxUMxa12_and_b1) );
  NOR2X1 U4096 ( .A(n221), .B(n4541), 
        .Y(output_p1_times_a1_mul_componentxUMxa14_and_b0) );
  NOR2X1 U4097 ( .A(n221), .B(n228), 
        .Y(output_p1_times_a1_mul_componentxUMxa3_and_b0) );
  NOR2X1 U4098 ( .A(n221), .B(n222), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b0) );
  NOR2X1 U4099 ( .A(n221), .B(n229), 
        .Y(output_p1_times_a1_mul_componentxUMxa2_and_b0) );
  NOR2X1 U4100 ( .A(n222), .B(n218), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b3) );
  NOR2X1 U4101 ( .A(n222), .B(n217), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b4) );
  NOR2X1 U4102 ( .A(n220), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b1) );
  NOR2X1 U4103 ( .A(n222), .B(n216), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b5) );
  NOR2X1 U4104 ( .A(n219), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b2) );
  NOR2X1 U4105 ( .A(n218), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b3) );
  NOR2X1 U4106 ( .A(n217), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b4) );
  NOR2X1 U4107 ( .A(n216), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b5) );
  NOR2X1 U4108 ( .A(n215), .B(n226), 
        .Y(output_p1_times_a1_mul_componentxUMxa5_and_b6) );
  NOR2X1 U4109 ( .A(n215), .B(n223), 
        .Y(output_p1_times_a1_mul_componentxUMxa8_and_b6) );
  NOR2X1 U4110 ( .A(n231), .B(n220), 
        .Y(output_p1_times_a1_mul_componentxUMxa0_and_b1) );
  NOR2X1 U4111 ( .A(n222), .B(n220), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b1) );
  NOR2X1 U4112 ( .A(n221), .B(n4545), 
        .Y(output_p1_times_a1_mul_componentxUMxa10_and_b0) );
  NOR2X1 U4113 ( .A(n221), .B(n4542), 
        .Y(output_p1_times_a1_mul_componentxUMxa13_and_b0) );
  NOR2X1 U4114 ( .A(n221), .B(n230), 
        .Y(output_p1_times_a1_mul_componentxUMxa1_and_b0) );
  XOR2X1 U4115 ( .A(n1338), .B(n1318), .Y(n4149) );
  XOR2X1 U4116 ( .A(n1336), .B(n1316), .Y(n4145) );
  XOR2X1 U4117 ( .A(n1230), .B(n1373), .Y(results_b0_b1_adderxn25) );
  XOR2X1 U4118 ( .A(n1334), .B(n1314), .Y(n4141) );
  XNOR2X1 U4119 ( .A(n1339), .B(n1319), .Y(n4151) );
  XNOR2X1 U4120 ( .A(n1337), .B(n1317), .Y(n4147) );
  XNOR2X1 U4121 ( .A(n1335), .B(n1315), .Y(n4143) );
  XOR2X1 U4122 ( .A(n1229), .B(n1372), .Y(results_b0_b1_adderxn22) );
  XOR2X1 U4123 ( .A(n1333), .B(n1313), .Y(n4138) );
  NOR2X1 U4124 ( .A(n231), .B(n221), 
        .Y(output_p1_times_a1_mul_componentxUMxfirst_vector[0]) );
  NOR2X1 U4125 ( .A(n216), .B(n4545), 
        .Y(output_p1_times_a1_mul_componentxUMxa10_and_b5) );
  NOR2X1 U4126 ( .A(n215), .B(n4545), 
        .Y(output_p1_times_a1_mul_componentxUMxa10_and_b6) );
  NOR2X1 U4127 ( .A(n218), .B(n4542), 
        .Y(output_p1_times_a1_mul_componentxUMxa13_and_b3) );
  NOR2X1 U4128 ( .A(n217), .B(n4544), 
        .Y(output_p1_times_a1_mul_componentxUMxa11_and_b4) );
  NOR2X1 U4129 ( .A(n216), .B(n4544), 
        .Y(output_p1_times_a1_mul_componentxUMxa11_and_b5) );
  NOR2X1 U4130 ( .A(n218), .B(n4543), 
        .Y(output_p1_times_a1_mul_componentxUMxa12_and_b3) );
  NOR2X1 U4131 ( .A(n217), .B(n4543), 
        .Y(output_p1_times_a1_mul_componentxUMxa12_and_b4) );
  NOR2X1 U4132 ( .A(n221), .B(n4540), 
        .Y(output_p1_times_a1_mul_componentxUMxa15_and_b0) );
  NOR2X1 U4133 ( .A(n220), .B(n4541), 
        .Y(output_p1_times_a1_mul_componentxUMxa14_and_b1) );
  NOR2X1 U4134 ( .A(n219), .B(n4541), 
        .Y(output_p1_times_a1_mul_componentxUMxa14_and_b2) );
  NOR2X1 U4135 ( .A(n220), .B(n4540), 
        .Y(output_p1_times_a1_mul_componentxUMxa15_and_b1) );
  NOR2X1 U4136 ( .A(n222), .B(n215), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b6) );
  NOR2X1 U4137 ( .A(n217), .B(n4542), 
        .Y(output_p1_times_a1_mul_componentxUMxa13_and_b4) );
  NOR2X1 U4138 ( .A(n221), .B(n4539), 
        .Y(output_p1_times_a1_mul_componentxUMxa16_and_b0) );
  XOR2X1 U4139 ( .A(output_p1_times_a1_mul_componentxUMxa14_and_b3), .B(n3185), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127715984_127849024_127850928)
         );
  NOR2X1 U4140 ( .A(n218), .B(n4541), 
        .Y(output_p1_times_a1_mul_componentxUMxa14_and_b3) );
  XOR2X1 U4141 ( .A(output_p1_times_a1_mul_componentxUMxa12_and_b5), 
        .B(output_p1_times_a1_mul_componentxUMxa13_and_b4), .Y(n3185) );
  NOR2X1 U4142 ( .A(n216), .B(n4543), 
        .Y(output_p1_times_a1_mul_componentxUMxa12_and_b5) );
  XOR2X1 U4143 ( .A(output_p1_times_a1_mul_componentxUMxa15_and_b2), 
        .B(output_p1_times_a1_mul_componentxUMxa16_and_b1), .Y(n3186) );
  NOR2X1 U4144 ( .A(n219), .B(n4540), 
        .Y(output_p1_times_a1_mul_componentxUMxa15_and_b2) );
  NOR2X1 U4145 ( .A(n220), .B(n4539), 
        .Y(output_p1_times_a1_mul_componentxUMxa16_and_b1) );
  XOR2X1 U4146 ( .A(output_p1_times_a1_mul_componentxUMxa11_and_b6), .B(n3184), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127636480_127638384_127714080)
         );
  NOR2X1 U4147 ( .A(n215), .B(n4544), 
        .Y(output_p1_times_a1_mul_componentxUMxa11_and_b6) );
  XOR2X1 U4148 ( .A(output_p1_times_a1_mul_componentxUMxa9_and_b8), 
        .B(output_p1_times_a1_mul_componentxUMxa10_and_b7), .Y(n3184) );
  NOR2X1 U4149 ( .A(n222), .B(n213), 
        .Y(output_p1_times_a1_mul_componentxUMxa9_and_b8) );
  XOR2X1 U4150 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127627616_127629520_127824000), 
        .B(n3246), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer2_128199816_128200040_128199984)
         );
  XOR2X1 U4151 ( .A(output_p1_times_a1_mul_componentxUMxa17_and_b0), .B(n3186), 
        .Y(output_p1_times_a1_mul_componentxUMxsum_layer1_127627616_127629520_127824000)
         );
  XOR2X1 U4152 ( 
        .A(output_p1_times_a1_mul_componentxUMxsum_layer1_127636480_127638384_127714080), 
        .B(output_p1_times_a1_mul_componentxUMxsum_layer1_127715984_127849024_127850928), 
        .Y(n3246) );
  NOR2X1 U4153 ( .A(n221), .B(n9), 
        .Y(output_p1_times_a1_mul_componentxUMxa17_and_b0) );
  NOR2X1 U4154 ( .A(n178), .B(n4439), 
        .Y(input_p1_times_b1_mul_componentxUMxa10_and_b1) );
  NOR2X1 U4155 ( .A(n199), .B(n4492), 
        .Y(input_p2_times_b2_mul_componentxUMxa10_and_b1) );
  NOR2X1 U4156 ( .A(n241), .B(n4598), 
        .Y(output_p2_times_a2_mul_componentxUMxa10_and_b1) );
  NOR2X1 U4157 ( .A(n269), .B(input_times_b0_mul_componentxn88), 
        .Y(input_times_b0_mul_componentxUMxa10_and_b1) );
  NOR2X1 U4158 ( .A(n179), .B(n4438), 
        .Y(input_p1_times_b1_mul_componentxUMxa11_and_b0) );
  NOR2X1 U4159 ( .A(n270), .B(input_times_b0_mul_componentxn87), 
        .Y(input_times_b0_mul_componentxUMxa11_and_b0) );
  NOR2X1 U4160 ( .A(n180), .B(n177), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b2) );
  NOR2X1 U4161 ( .A(n201), .B(n198), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b2) );
  NOR2X1 U4162 ( .A(n243), .B(n240), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b2) );
  NOR2X1 U4163 ( .A(n271), .B(n268), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b2) );
  NOR2X1 U4164 ( .A(n177), .B(n4439), 
        .Y(input_p1_times_b1_mul_componentxUMxa10_and_b2) );
  NOR2X1 U4165 ( .A(n198), .B(n4492), 
        .Y(input_p2_times_b2_mul_componentxUMxa10_and_b2) );
  NOR2X1 U4166 ( .A(n240), .B(n4598), 
        .Y(output_p2_times_a2_mul_componentxUMxa10_and_b2) );
  NOR2X1 U4167 ( .A(n268), .B(input_times_b0_mul_componentxn88), 
        .Y(input_times_b0_mul_componentxUMxa10_and_b2) );
  NOR2X1 U4168 ( .A(n176), .B(n4439), 
        .Y(input_p1_times_b1_mul_componentxUMxa10_and_b3) );
  NOR2X1 U4169 ( .A(n197), .B(n4492), 
        .Y(input_p2_times_b2_mul_componentxUMxa10_and_b3) );
  NOR2X1 U4170 ( .A(n239), .B(n4598), 
        .Y(output_p2_times_a2_mul_componentxUMxa10_and_b3) );
  NOR2X1 U4171 ( .A(n267), .B(input_times_b0_mul_componentxn88), 
        .Y(input_times_b0_mul_componentxUMxa10_and_b3) );
  NOR2X1 U4172 ( .A(n175), .B(n4439), 
        .Y(input_p1_times_b1_mul_componentxUMxa10_and_b4) );
  NOR2X1 U4173 ( .A(n196), .B(n4492), 
        .Y(input_p2_times_b2_mul_componentxUMxa10_and_b4) );
  NOR2X1 U4174 ( .A(n238), .B(n4598), 
        .Y(output_p2_times_a2_mul_componentxUMxa10_and_b4) );
  NOR2X1 U4175 ( .A(n266), .B(input_times_b0_mul_componentxn88), 
        .Y(input_times_b0_mul_componentxUMxa10_and_b4) );
  NOR2X1 U4176 ( .A(n178), .B(n4436), 
        .Y(input_p1_times_b1_mul_componentxUMxa13_and_b1) );
  NOR2X1 U4177 ( .A(n269), .B(input_times_b0_mul_componentxn85), 
        .Y(input_times_b0_mul_componentxUMxa13_and_b1) );
  NOR2X1 U4178 ( .A(n177), .B(n4436), 
        .Y(input_p1_times_b1_mul_componentxUMxa13_and_b2) );
  NOR2X1 U4179 ( .A(n268), .B(input_times_b0_mul_componentxn85), 
        .Y(input_times_b0_mul_componentxUMxa13_and_b2) );
  NOR2X1 U4180 ( .A(n199), .B(n4489), 
        .Y(input_p2_times_b2_mul_componentxUMxa13_and_b1) );
  NOR2X1 U4181 ( .A(n241), .B(n4595), 
        .Y(output_p2_times_a2_mul_componentxUMxa13_and_b1) );
  NOR2X1 U4182 ( .A(n198), .B(n4489), 
        .Y(input_p2_times_b2_mul_componentxUMxa13_and_b2) );
  NOR2X1 U4183 ( .A(n240), .B(n4595), 
        .Y(output_p2_times_a2_mul_componentxUMxa13_and_b2) );
  NOR2X1 U4184 ( .A(n178), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b1) );
  NOR2X1 U4185 ( .A(n199), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b1) );
  NOR2X1 U4186 ( .A(n241), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b1) );
  NOR2X1 U4187 ( .A(n269), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b1) );
  NOR2X1 U4188 ( .A(n178), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b1) );
  NOR2X1 U4189 ( .A(n199), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b1) );
  NOR2X1 U4190 ( .A(n241), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b1) );
  NOR2X1 U4191 ( .A(n269), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b1) );
  NOR2X1 U4192 ( .A(n177), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b2) );
  NOR2X1 U4193 ( .A(n198), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b2) );
  NOR2X1 U4194 ( .A(n240), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b2) );
  NOR2X1 U4195 ( .A(n268), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b2) );
  NOR2X1 U4196 ( .A(n177), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b2) );
  NOR2X1 U4197 ( .A(n198), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b2) );
  NOR2X1 U4198 ( .A(n240), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b2) );
  NOR2X1 U4199 ( .A(n268), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b2) );
  NOR2X1 U4200 ( .A(n177), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b2) );
  NOR2X1 U4201 ( .A(n198), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b2) );
  NOR2X1 U4202 ( .A(n240), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b2) );
  NOR2X1 U4203 ( .A(n268), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b2) );
  NOR2X1 U4204 ( .A(n176), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b3) );
  NOR2X1 U4205 ( .A(n197), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b3) );
  NOR2X1 U4206 ( .A(n239), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b3) );
  NOR2X1 U4207 ( .A(n267), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b3) );
  NOR2X1 U4208 ( .A(n176), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b3) );
  NOR2X1 U4209 ( .A(n197), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b3) );
  NOR2X1 U4210 ( .A(n239), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b3) );
  NOR2X1 U4211 ( .A(n267), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b3) );
  NOR2X1 U4212 ( .A(n176), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b3) );
  NOR2X1 U4213 ( .A(n197), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b3) );
  NOR2X1 U4214 ( .A(n239), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b3) );
  NOR2X1 U4215 ( .A(n267), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b3) );
  NOR2X1 U4216 ( .A(n175), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b4) );
  NOR2X1 U4217 ( .A(n196), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b4) );
  NOR2X1 U4218 ( .A(n238), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b4) );
  NOR2X1 U4219 ( .A(n266), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b4) );
  NOR2X1 U4220 ( .A(n175), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b4) );
  NOR2X1 U4221 ( .A(n196), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b4) );
  NOR2X1 U4222 ( .A(n238), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b4) );
  NOR2X1 U4223 ( .A(n266), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b4) );
  NOR2X1 U4224 ( .A(n175), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b4) );
  NOR2X1 U4225 ( .A(n196), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b4) );
  NOR2X1 U4226 ( .A(n238), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b4) );
  NOR2X1 U4227 ( .A(n266), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b4) );
  NOR2X1 U4228 ( .A(n174), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b5) );
  NOR2X1 U4229 ( .A(n195), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b5) );
  NOR2X1 U4230 ( .A(n237), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b5) );
  NOR2X1 U4231 ( .A(n265), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b5) );
  NOR2X1 U4232 ( .A(n174), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b5) );
  NOR2X1 U4233 ( .A(n195), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b5) );
  NOR2X1 U4234 ( .A(n237), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b5) );
  NOR2X1 U4235 ( .A(n265), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b5) );
  NOR2X1 U4236 ( .A(n174), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b5) );
  NOR2X1 U4237 ( .A(n195), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b5) );
  NOR2X1 U4238 ( .A(n237), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b5) );
  NOR2X1 U4239 ( .A(n265), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b5) );
  NOR2X1 U4240 ( .A(n172), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b7) );
  NOR2X1 U4241 ( .A(n173), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b6) );
  NOR2X1 U4242 ( .A(n194), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b6) );
  NOR2X1 U4243 ( .A(n236), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b6) );
  NOR2X1 U4244 ( .A(n263), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b7) );
  NOR2X1 U4245 ( .A(n264), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b6) );
  NOR2X1 U4246 ( .A(n173), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b6) );
  NOR2X1 U4247 ( .A(n194), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b6) );
  NOR2X1 U4248 ( .A(n236), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b6) );
  NOR2X1 U4249 ( .A(n264), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b6) );
  NOR2X1 U4250 ( .A(n193), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b7) );
  NOR2X1 U4251 ( .A(n235), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b7) );
  NOR2X1 U4252 ( .A(n172), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b7) );
  NOR2X1 U4253 ( .A(n263), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b7) );
  NOR2X1 U4254 ( .A(n178), .B(n4438), 
        .Y(input_p1_times_b1_mul_componentxUMxa11_and_b1) );
  NOR2X1 U4255 ( .A(n269), .B(input_times_b0_mul_componentxn87), 
        .Y(input_times_b0_mul_componentxUMxa11_and_b1) );
  NOR2X1 U4256 ( .A(n177), .B(n4438), 
        .Y(input_p1_times_b1_mul_componentxUMxa11_and_b2) );
  NOR2X1 U4257 ( .A(n268), .B(input_times_b0_mul_componentxn87), 
        .Y(input_times_b0_mul_componentxUMxa11_and_b2) );
  NOR2X1 U4258 ( .A(n176), .B(n4438), 
        .Y(input_p1_times_b1_mul_componentxUMxa11_and_b3) );
  NOR2X1 U4259 ( .A(n267), .B(input_times_b0_mul_componentxn87), 
        .Y(input_times_b0_mul_componentxUMxa11_and_b3) );
  NOR2X1 U4260 ( .A(n179), .B(n4437), 
        .Y(input_p1_times_b1_mul_componentxUMxa12_and_b0) );
  NOR2X1 U4261 ( .A(n270), .B(input_times_b0_mul_componentxn86), 
        .Y(input_times_b0_mul_componentxUMxa12_and_b0) );
  NOR2X1 U4262 ( .A(n177), .B(n4437), 
        .Y(input_p1_times_b1_mul_componentxUMxa12_and_b2) );
  NOR2X1 U4263 ( .A(n268), .B(input_times_b0_mul_componentxn86), 
        .Y(input_times_b0_mul_componentxUMxa12_and_b2) );
  NOR2X1 U4264 ( .A(n200), .B(n4491), 
        .Y(input_p2_times_b2_mul_componentxUMxa11_and_b0) );
  NOR2X1 U4265 ( .A(n242), .B(n4597), 
        .Y(output_p2_times_a2_mul_componentxUMxa11_and_b0) );
  NOR2X1 U4266 ( .A(n199), .B(n4491), 
        .Y(input_p2_times_b2_mul_componentxUMxa11_and_b1) );
  NOR2X1 U4267 ( .A(n241), .B(n4597), 
        .Y(output_p2_times_a2_mul_componentxUMxa11_and_b1) );
  NOR2X1 U4268 ( .A(n198), .B(n4491), 
        .Y(input_p2_times_b2_mul_componentxUMxa11_and_b2) );
  NOR2X1 U4269 ( .A(n240), .B(n4597), 
        .Y(output_p2_times_a2_mul_componentxUMxa11_and_b2) );
  NOR2X1 U4270 ( .A(n197), .B(n4491), 
        .Y(input_p2_times_b2_mul_componentxUMxa11_and_b3) );
  NOR2X1 U4271 ( .A(n239), .B(n4597), 
        .Y(output_p2_times_a2_mul_componentxUMxa11_and_b3) );
  NOR2X1 U4272 ( .A(n200), .B(n4490), 
        .Y(input_p2_times_b2_mul_componentxUMxa12_and_b0) );
  NOR2X1 U4273 ( .A(n242), .B(n4596), 
        .Y(output_p2_times_a2_mul_componentxUMxa12_and_b0) );
  NOR2X1 U4274 ( .A(n198), .B(n4490), 
        .Y(input_p2_times_b2_mul_componentxUMxa12_and_b2) );
  NOR2X1 U4275 ( .A(n240), .B(n4596), 
        .Y(output_p2_times_a2_mul_componentxUMxa12_and_b2) );
  NOR2X1 U4276 ( .A(n179), .B(n4434), 
        .Y(input_p1_times_b1_mul_componentxUMxa15_and_b0) );
  NOR2X1 U4277 ( .A(n270), .B(input_times_b0_mul_componentxn83), 
        .Y(input_times_b0_mul_componentxUMxa15_and_b0) );
  NOR2X1 U4278 ( .A(n179), .B(n4435), 
        .Y(input_p1_times_b1_mul_componentxUMxa14_and_b0) );
  NOR2X1 U4279 ( .A(n270), .B(input_times_b0_mul_componentxn84), 
        .Y(input_times_b0_mul_componentxUMxa14_and_b0) );
  NOR2X1 U4280 ( .A(n178), .B(n4437), 
        .Y(input_p1_times_b1_mul_componentxUMxa12_and_b1) );
  NOR2X1 U4281 ( .A(n269), .B(input_times_b0_mul_componentxn86), 
        .Y(input_times_b0_mul_componentxUMxa12_and_b1) );
  NOR2X1 U4282 ( .A(n200), .B(n4487), 
        .Y(input_p2_times_b2_mul_componentxUMxa15_and_b0) );
  NOR2X1 U4283 ( .A(n242), .B(n4593), 
        .Y(output_p2_times_a2_mul_componentxUMxa15_and_b0) );
  NOR2X1 U4284 ( .A(n199), .B(n4490), 
        .Y(input_p2_times_b2_mul_componentxUMxa12_and_b1) );
  NOR2X1 U4285 ( .A(n241), .B(n4596), 
        .Y(output_p2_times_a2_mul_componentxUMxa12_and_b1) );
  NOR2X1 U4286 ( .A(n200), .B(n4488), 
        .Y(input_p2_times_b2_mul_componentxUMxa14_and_b0) );
  NOR2X1 U4287 ( .A(n242), .B(n4594), 
        .Y(output_p2_times_a2_mul_componentxUMxa14_and_b0) );
  NOR2X1 U4288 ( .A(n189), .B(n175), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b4) );
  NOR2X1 U4289 ( .A(n280), .B(n266), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b4) );
  NOR2X1 U4290 ( .A(n189), .B(n174), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b5) );
  NOR2X1 U4291 ( .A(n280), .B(n265), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b5) );
  NOR2X1 U4292 ( .A(n189), .B(n176), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b3) );
  NOR2X1 U4293 ( .A(n280), .B(n267), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b3) );
  NOR2X1 U4294 ( .A(n189), .B(n171), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b8) );
  NOR2X1 U4295 ( .A(n189), .B(n172), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b7) );
  NOR2X1 U4296 ( .A(n280), .B(n262), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b8) );
  NOR2X1 U4297 ( .A(n280), .B(n263), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b7) );
  NOR2X1 U4298 ( .A(n189), .B(n173), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b6) );
  NOR2X1 U4299 ( .A(n280), .B(n264), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b6) );
  NOR2X1 U4300 ( .A(n210), .B(n196), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b4) );
  NOR2X1 U4301 ( .A(n252), .B(n238), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b4) );
  NOR2X1 U4302 ( .A(n210), .B(n195), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b5) );
  NOR2X1 U4303 ( .A(n252), .B(n237), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b5) );
  NOR2X1 U4304 ( .A(n210), .B(n197), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b3) );
  NOR2X1 U4305 ( .A(n252), .B(n239), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b3) );
  NOR2X1 U4306 ( .A(n210), .B(n192), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b8) );
  NOR2X1 U4307 ( .A(n210), .B(n193), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b7) );
  NOR2X1 U4308 ( .A(n252), .B(n234), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b8) );
  NOR2X1 U4309 ( .A(n252), .B(n235), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b7) );
  NOR2X1 U4310 ( .A(n210), .B(n194), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b6) );
  NOR2X1 U4311 ( .A(n252), .B(n236), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b6) );
  NOR2X1 U4312 ( .A(n179), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b0) );
  NOR2X1 U4313 ( .A(n200), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b0) );
  NOR2X1 U4314 ( .A(n242), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b0) );
  NOR2X1 U4315 ( .A(n270), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b0) );
  NOR2X1 U4316 ( .A(n179), .B(n180), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b0) );
  NOR2X1 U4317 ( .A(n200), .B(n201), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b0) );
  NOR2X1 U4318 ( .A(n242), .B(n243), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b0) );
  NOR2X1 U4319 ( .A(n270), .B(n271), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b0) );
  NOR2X1 U4320 ( .A(n177), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b2) );
  NOR2X1 U4321 ( .A(n198), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b2) );
  NOR2X1 U4322 ( .A(n240), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b2) );
  NOR2X1 U4323 ( .A(n268), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b2) );
  NOR2X1 U4324 ( .A(n177), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b2) );
  NOR2X1 U4325 ( .A(n198), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b2) );
  NOR2X1 U4326 ( .A(n240), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b2) );
  NOR2X1 U4327 ( .A(n268), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b2) );
  NOR2X1 U4328 ( .A(n176), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b3) );
  NOR2X1 U4329 ( .A(n197), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b3) );
  NOR2X1 U4330 ( .A(n239), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b3) );
  NOR2X1 U4331 ( .A(n267), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b3) );
  NOR2X1 U4332 ( .A(n176), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b3) );
  NOR2X1 U4333 ( .A(n197), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b3) );
  NOR2X1 U4334 ( .A(n239), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b3) );
  NOR2X1 U4335 ( .A(n267), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b3) );
  NOR2X1 U4336 ( .A(n175), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b4) );
  NOR2X1 U4337 ( .A(n196), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b4) );
  NOR2X1 U4338 ( .A(n238), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b4) );
  NOR2X1 U4339 ( .A(n266), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b4) );
  NOR2X1 U4340 ( .A(n175), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b4) );
  NOR2X1 U4341 ( .A(n196), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b4) );
  NOR2X1 U4342 ( .A(n238), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b4) );
  NOR2X1 U4343 ( .A(n266), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b4) );
  NOR2X1 U4344 ( .A(n174), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b5) );
  NOR2X1 U4345 ( .A(n195), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b5) );
  NOR2X1 U4346 ( .A(n237), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b5) );
  NOR2X1 U4347 ( .A(n265), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b5) );
  NOR2X1 U4348 ( .A(n174), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b5) );
  NOR2X1 U4349 ( .A(n195), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b5) );
  NOR2X1 U4350 ( .A(n237), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b5) );
  NOR2X1 U4351 ( .A(n265), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b5) );
  NOR2X1 U4352 ( .A(n173), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b6) );
  NOR2X1 U4353 ( .A(n264), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b6) );
  NOR2X1 U4354 ( .A(n173), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b6) );
  NOR2X1 U4355 ( .A(n194), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b6) );
  NOR2X1 U4356 ( .A(n236), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b6) );
  NOR2X1 U4357 ( .A(n264), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b6) );
  NOR2X1 U4358 ( .A(n179), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b0) );
  NOR2X1 U4359 ( .A(n200), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b0) );
  NOR2X1 U4360 ( .A(n242), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b0) );
  NOR2X1 U4361 ( .A(n270), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b0) );
  NOR2X1 U4362 ( .A(n179), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b0) );
  NOR2X1 U4363 ( .A(n200), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b0) );
  NOR2X1 U4364 ( .A(n242), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b0) );
  NOR2X1 U4365 ( .A(n270), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b0) );
  NOR2X1 U4366 ( .A(n180), .B(n176), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b3) );
  NOR2X1 U4367 ( .A(n201), .B(n197), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b3) );
  NOR2X1 U4368 ( .A(n243), .B(n239), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b3) );
  NOR2X1 U4369 ( .A(n271), .B(n267), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b3) );
  NOR2X1 U4370 ( .A(n172), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b7) );
  NOR2X1 U4371 ( .A(n193), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b7) );
  NOR2X1 U4372 ( .A(n235), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b7) );
  NOR2X1 U4373 ( .A(n263), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b7) );
  NOR2X1 U4374 ( .A(n180), .B(n175), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b4) );
  NOR2X1 U4375 ( .A(n201), .B(n196), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b4) );
  NOR2X1 U4376 ( .A(n243), .B(n238), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b4) );
  NOR2X1 U4377 ( .A(n271), .B(n266), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b4) );
  NOR2X1 U4378 ( .A(n178), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b1) );
  NOR2X1 U4379 ( .A(n199), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b1) );
  NOR2X1 U4380 ( .A(n241), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b1) );
  NOR2X1 U4381 ( .A(n269), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b1) );
  NOR2X1 U4382 ( .A(n178), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b1) );
  NOR2X1 U4383 ( .A(n199), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b1) );
  NOR2X1 U4384 ( .A(n241), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b1) );
  NOR2X1 U4385 ( .A(n269), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b1) );
  NOR2X1 U4386 ( .A(n180), .B(n174), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b5) );
  NOR2X1 U4387 ( .A(n201), .B(n195), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b5) );
  NOR2X1 U4388 ( .A(n243), .B(n237), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b5) );
  NOR2X1 U4389 ( .A(n271), .B(n265), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b5) );
  NOR2X1 U4390 ( .A(n177), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b2) );
  NOR2X1 U4391 ( .A(n198), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b2) );
  NOR2X1 U4392 ( .A(n240), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b2) );
  NOR2X1 U4393 ( .A(n268), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b2) );
  NOR2X1 U4394 ( .A(n177), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b2) );
  NOR2X1 U4395 ( .A(n198), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b2) );
  NOR2X1 U4396 ( .A(n240), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b2) );
  NOR2X1 U4397 ( .A(n268), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b2) );
  NOR2X1 U4398 ( .A(n177), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b2) );
  NOR2X1 U4399 ( .A(n198), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b2) );
  NOR2X1 U4400 ( .A(n240), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b2) );
  NOR2X1 U4401 ( .A(n268), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b2) );
  NOR2X1 U4402 ( .A(n176), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b3) );
  NOR2X1 U4403 ( .A(n197), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b3) );
  NOR2X1 U4404 ( .A(n239), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b3) );
  NOR2X1 U4405 ( .A(n267), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b3) );
  NOR2X1 U4406 ( .A(n176), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b3) );
  NOR2X1 U4407 ( .A(n197), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b3) );
  NOR2X1 U4408 ( .A(n239), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b3) );
  NOR2X1 U4409 ( .A(n267), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b3) );
  NOR2X1 U4410 ( .A(n176), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b3) );
  NOR2X1 U4411 ( .A(n197), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b3) );
  NOR2X1 U4412 ( .A(n239), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b3) );
  NOR2X1 U4413 ( .A(n267), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b3) );
  NOR2X1 U4414 ( .A(n175), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b4) );
  NOR2X1 U4415 ( .A(n196), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b4) );
  NOR2X1 U4416 ( .A(n238), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b4) );
  NOR2X1 U4417 ( .A(n266), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b4) );
  NOR2X1 U4418 ( .A(n175), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b4) );
  NOR2X1 U4419 ( .A(n196), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b4) );
  NOR2X1 U4420 ( .A(n238), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b4) );
  NOR2X1 U4421 ( .A(n266), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b4) );
  NOR2X1 U4422 ( .A(n174), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b5) );
  NOR2X1 U4423 ( .A(n195), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b5) );
  NOR2X1 U4424 ( .A(n237), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b5) );
  NOR2X1 U4425 ( .A(n265), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b5) );
  NOR2X1 U4426 ( .A(n174), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b5) );
  NOR2X1 U4427 ( .A(n265), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b5) );
  NOR2X1 U4428 ( .A(n178), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b1) );
  NOR2X1 U4429 ( .A(n199), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b1) );
  NOR2X1 U4430 ( .A(n241), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b1) );
  NOR2X1 U4431 ( .A(n269), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b1) );
  NOR2X1 U4432 ( .A(n178), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b1) );
  NOR2X1 U4433 ( .A(n199), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b1) );
  NOR2X1 U4434 ( .A(n241), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b1) );
  NOR2X1 U4435 ( .A(n269), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b1) );
  NOR2X1 U4436 ( .A(n180), .B(n178), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b1) );
  NOR2X1 U4437 ( .A(n201), .B(n199), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b1) );
  NOR2X1 U4438 ( .A(n243), .B(n241), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b1) );
  NOR2X1 U4439 ( .A(n271), .B(n269), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b1) );
  NOR2X1 U4440 ( .A(n179), .B(n4439), 
        .Y(input_p1_times_b1_mul_componentxUMxa10_and_b0) );
  NOR2X1 U4441 ( .A(n200), .B(n4492), 
        .Y(input_p2_times_b2_mul_componentxUMxa10_and_b0) );
  NOR2X1 U4442 ( .A(n242), .B(n4598), 
        .Y(output_p2_times_a2_mul_componentxUMxa10_and_b0) );
  NOR2X1 U4443 ( .A(n270), .B(input_times_b0_mul_componentxn88), 
        .Y(input_times_b0_mul_componentxUMxa10_and_b0) );
  NOR2X1 U4444 ( .A(n179), .B(n4436), 
        .Y(input_p1_times_b1_mul_componentxUMxa13_and_b0) );
  NOR2X1 U4445 ( .A(n270), .B(input_times_b0_mul_componentxn85), 
        .Y(input_times_b0_mul_componentxUMxa13_and_b0) );
  NOR2X1 U4446 ( .A(n200), .B(n4489), 
        .Y(input_p2_times_b2_mul_componentxUMxa13_and_b0) );
  NOR2X1 U4447 ( .A(n242), .B(n4595), 
        .Y(output_p2_times_a2_mul_componentxUMxa13_and_b0) );
  NOR2X1 U4448 ( .A(n179), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b0) );
  NOR2X1 U4449 ( .A(n200), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b0) );
  NOR2X1 U4450 ( .A(n242), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b0) );
  NOR2X1 U4451 ( .A(n270), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b0) );
  NOR2X1 U4452 ( .A(n179), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b0) );
  NOR2X1 U4453 ( .A(n200), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b0) );
  NOR2X1 U4454 ( .A(n242), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b0) );
  NOR2X1 U4455 ( .A(n270), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b0) );
  NOR2X1 U4456 ( .A(n4422), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b10) );
  NOR2X1 U4457 ( .A(n4475), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b10) );
  NOR2X1 U4458 ( .A(n4581), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b10) );
  NOR2X1 U4459 ( .A(input_times_b0_mul_componentxn71), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b10) );
  NOR2X1 U4460 ( .A(n4422), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b10) );
  NOR2X1 U4461 ( .A(n4475), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b10) );
  NOR2X1 U4462 ( .A(n4581), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b10) );
  NOR2X1 U4463 ( .A(input_times_b0_mul_componentxn71), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b10) );
  NOR2X1 U4464 ( .A(n174), .B(n4439), 
        .Y(input_p1_times_b1_mul_componentxUMxa10_and_b5) );
  NOR2X1 U4465 ( .A(n195), .B(n4492), 
        .Y(input_p2_times_b2_mul_componentxUMxa10_and_b5) );
  NOR2X1 U4466 ( .A(n237), .B(n4598), 
        .Y(output_p2_times_a2_mul_componentxUMxa10_and_b5) );
  NOR2X1 U4467 ( .A(n265), .B(input_times_b0_mul_componentxn88), 
        .Y(input_times_b0_mul_componentxUMxa10_and_b5) );
  NOR2X1 U4468 ( .A(n173), .B(n4439), 
        .Y(input_p1_times_b1_mul_componentxUMxa10_and_b6) );
  NOR2X1 U4469 ( .A(n194), .B(n4492), 
        .Y(input_p2_times_b2_mul_componentxUMxa10_and_b6) );
  NOR2X1 U4470 ( .A(n236), .B(n4598), 
        .Y(output_p2_times_a2_mul_componentxUMxa10_and_b6) );
  NOR2X1 U4471 ( .A(n264), .B(input_times_b0_mul_componentxn88), 
        .Y(input_times_b0_mul_componentxUMxa10_and_b6) );
  NOR2X1 U4472 ( .A(n4421), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b11) );
  NOR2X1 U4473 ( .A(n4474), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b11) );
  NOR2X1 U4474 ( .A(n4580), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b11) );
  NOR2X1 U4475 ( .A(input_times_b0_mul_componentxn70), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b11) );
  NOR2X1 U4476 ( .A(n4420), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b12) );
  NOR2X1 U4477 ( .A(n4473), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b12) );
  NOR2X1 U4478 ( .A(n4579), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b12) );
  NOR2X1 U4479 ( .A(input_times_b0_mul_componentxn69), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b12) );
  NOR2X1 U4480 ( .A(n176), .B(n4436), 
        .Y(input_p1_times_b1_mul_componentxUMxa13_and_b3) );
  NOR2X1 U4481 ( .A(n267), .B(input_times_b0_mul_componentxn85), 
        .Y(input_times_b0_mul_componentxUMxa13_and_b3) );
  NOR2X1 U4482 ( .A(n197), .B(n4489), 
        .Y(input_p2_times_b2_mul_componentxUMxa13_and_b3) );
  NOR2X1 U4483 ( .A(n239), .B(n4595), 
        .Y(output_p2_times_a2_mul_componentxUMxa13_and_b3) );
  NOR2X1 U4484 ( .A(n178), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b1) );
  NOR2X1 U4485 ( .A(n199), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b1) );
  NOR2X1 U4486 ( .A(n241), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b1) );
  NOR2X1 U4487 ( .A(n269), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b1) );
  NOR2X1 U4488 ( .A(n171), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b8) );
  NOR2X1 U4489 ( .A(n262), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b8) );
  NOR2X1 U4490 ( .A(n170), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b9) );
  NOR2X1 U4491 ( .A(n261), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b9) );
  NOR2X1 U4492 ( .A(n173), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b6) );
  NOR2X1 U4493 ( .A(n194), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b6) );
  NOR2X1 U4494 ( .A(n236), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b6) );
  NOR2X1 U4495 ( .A(n264), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b6) );
  NOR2X1 U4496 ( .A(n192), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b8) );
  NOR2X1 U4497 ( .A(n234), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b8) );
  NOR2X1 U4498 ( .A(n191), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b9) );
  NOR2X1 U4499 ( .A(n233), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b9) );
  NOR2X1 U4500 ( .A(n172), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b7) );
  NOR2X1 U4501 ( .A(n193), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b7) );
  NOR2X1 U4502 ( .A(n235), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b7) );
  NOR2X1 U4503 ( .A(n263), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b7) );
  NOR2X1 U4504 ( .A(n193), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b7) );
  NOR2X1 U4505 ( .A(n235), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b7) );
  NOR2X1 U4506 ( .A(n171), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b8) );
  NOR2X1 U4507 ( .A(n262), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b8) );
  NOR2X1 U4508 ( .A(n170), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b9) );
  NOR2X1 U4509 ( .A(n261), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b9) );
  NOR2X1 U4510 ( .A(n192), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b8) );
  NOR2X1 U4511 ( .A(n234), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b8) );
  NOR2X1 U4512 ( .A(n191), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b9) );
  NOR2X1 U4513 ( .A(n233), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b9) );
  NOR2X1 U4514 ( .A(n171), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b8) );
  NOR2X1 U4515 ( .A(n262), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b8) );
  NOR2X1 U4516 ( .A(n4422), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b10) );
  NOR2X1 U4517 ( .A(n4475), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b10) );
  NOR2X1 U4518 ( .A(n4581), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b10) );
  NOR2X1 U4519 ( .A(input_times_b0_mul_componentxn71), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b10) );
  NOR2X1 U4520 ( .A(n189), .B(n4422), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b10) );
  NOR2X1 U4521 ( .A(n210), .B(n4475), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b10) );
  NOR2X1 U4522 ( .A(n252), .B(n4581), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b10) );
  NOR2X1 U4523 ( .A(n280), .B(input_times_b0_mul_componentxn71), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b10) );
  NOR2X1 U4524 ( .A(n4422), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b10) );
  NOR2X1 U4525 ( .A(n4475), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b10) );
  NOR2X1 U4526 ( .A(n4581), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b10) );
  NOR2X1 U4527 ( .A(input_times_b0_mul_componentxn71), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b10) );
  NOR2X1 U4528 ( .A(n4421), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b11) );
  NOR2X1 U4529 ( .A(n4474), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b11) );
  NOR2X1 U4530 ( .A(n4580), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b11) );
  NOR2X1 U4531 ( .A(input_times_b0_mul_componentxn70), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b11) );
  NOR2X1 U4532 ( .A(n189), .B(n4421), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b11) );
  NOR2X1 U4533 ( .A(n210), .B(n4474), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b11) );
  NOR2X1 U4534 ( .A(n252), .B(n4580), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b11) );
  NOR2X1 U4535 ( .A(n280), .B(input_times_b0_mul_componentxn70), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b11) );
  NOR2X1 U4536 ( .A(n4421), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b11) );
  NOR2X1 U4537 ( .A(n4474), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b11) );
  NOR2X1 U4538 ( .A(n4580), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b11) );
  NOR2X1 U4539 ( .A(input_times_b0_mul_componentxn70), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b11) );
  NOR2X1 U4540 ( .A(n175), .B(n4438), 
        .Y(input_p1_times_b1_mul_componentxUMxa11_and_b4) );
  NOR2X1 U4541 ( .A(n266), .B(input_times_b0_mul_componentxn87), 
        .Y(input_times_b0_mul_componentxUMxa11_and_b4) );
  NOR2X1 U4542 ( .A(n174), .B(n4438), 
        .Y(input_p1_times_b1_mul_componentxUMxa11_and_b5) );
  NOR2X1 U4543 ( .A(n265), .B(input_times_b0_mul_componentxn87), 
        .Y(input_times_b0_mul_componentxUMxa11_and_b5) );
  NOR2X1 U4544 ( .A(n176), .B(n4437), 
        .Y(input_p1_times_b1_mul_componentxUMxa12_and_b3) );
  NOR2X1 U4545 ( .A(n267), .B(input_times_b0_mul_componentxn86), 
        .Y(input_times_b0_mul_componentxUMxa12_and_b3) );
  NOR2X1 U4546 ( .A(n175), .B(n4437), 
        .Y(input_p1_times_b1_mul_componentxUMxa12_and_b4) );
  NOR2X1 U4547 ( .A(n266), .B(input_times_b0_mul_componentxn86), 
        .Y(input_times_b0_mul_componentxUMxa12_and_b4) );
  NOR2X1 U4548 ( .A(n189), .B(n4420), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b12) );
  NOR2X1 U4549 ( .A(n210), .B(n4473), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b12) );
  NOR2X1 U4550 ( .A(n252), .B(n4579), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b12) );
  NOR2X1 U4551 ( .A(n280), .B(input_times_b0_mul_componentxn69), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b12) );
  NOR2X1 U4552 ( .A(n196), .B(n4491), 
        .Y(input_p2_times_b2_mul_componentxUMxa11_and_b4) );
  NOR2X1 U4553 ( .A(n238), .B(n4597), 
        .Y(output_p2_times_a2_mul_componentxUMxa11_and_b4) );
  NOR2X1 U4554 ( .A(n195), .B(n4491), 
        .Y(input_p2_times_b2_mul_componentxUMxa11_and_b5) );
  NOR2X1 U4555 ( .A(n237), .B(n4597), 
        .Y(output_p2_times_a2_mul_componentxUMxa11_and_b5) );
  NOR2X1 U4556 ( .A(n197), .B(n4490), 
        .Y(input_p2_times_b2_mul_componentxUMxa12_and_b3) );
  NOR2X1 U4557 ( .A(n239), .B(n4596), 
        .Y(output_p2_times_a2_mul_componentxUMxa12_and_b3) );
  NOR2X1 U4558 ( .A(n196), .B(n4490), 
        .Y(input_p2_times_b2_mul_componentxUMxa12_and_b4) );
  NOR2X1 U4559 ( .A(n238), .B(n4596), 
        .Y(output_p2_times_a2_mul_componentxUMxa12_and_b4) );
  NOR2X1 U4560 ( .A(n280), .B(input_times_b0_mul_componentxn68), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b13) );
  NOR2X1 U4561 ( .A(n189), .B(n4419), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b13) );
  NOR2X1 U4562 ( .A(n210), .B(n4472), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b13) );
  NOR2X1 U4563 ( .A(n252), .B(n4578), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b13) );
  NOR2X1 U4564 ( .A(n178), .B(n4435), 
        .Y(input_p1_times_b1_mul_componentxUMxa14_and_b1) );
  NOR2X1 U4565 ( .A(n269), .B(input_times_b0_mul_componentxn84), 
        .Y(input_times_b0_mul_componentxUMxa14_and_b1) );
  NOR2X1 U4566 ( .A(n177), .B(n4435), 
        .Y(input_p1_times_b1_mul_componentxUMxa14_and_b2) );
  NOR2X1 U4567 ( .A(n268), .B(input_times_b0_mul_componentxn84), 
        .Y(input_times_b0_mul_componentxUMxa14_and_b2) );
  NOR2X1 U4568 ( .A(n199), .B(n4488), 
        .Y(input_p2_times_b2_mul_componentxUMxa14_and_b1) );
  NOR2X1 U4569 ( .A(n241), .B(n4594), 
        .Y(output_p2_times_a2_mul_componentxUMxa14_and_b1) );
  NOR2X1 U4570 ( .A(n198), .B(n4488), 
        .Y(input_p2_times_b2_mul_componentxUMxa14_and_b2) );
  NOR2X1 U4571 ( .A(n240), .B(n4594), 
        .Y(output_p2_times_a2_mul_componentxUMxa14_and_b2) );
  NOR2X1 U4572 ( .A(n178), .B(n4434), 
        .Y(input_p1_times_b1_mul_componentxUMxa15_and_b1) );
  NOR2X1 U4573 ( .A(n269), .B(input_times_b0_mul_componentxn83), 
        .Y(input_times_b0_mul_componentxUMxa15_and_b1) );
  NOR2X1 U4574 ( .A(n189), .B(n177), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b2) );
  NOR2X1 U4575 ( .A(n280), .B(n268), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b2) );
  NOR2X1 U4576 ( .A(n189), .B(n170), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b9) );
  NOR2X1 U4577 ( .A(n280), .B(n261), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b9) );
  NOR2X1 U4578 ( .A(n210), .B(n198), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b2) );
  NOR2X1 U4579 ( .A(n252), .B(n240), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b2) );
  NOR2X1 U4580 ( .A(n210), .B(n191), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b9) );
  NOR2X1 U4581 ( .A(n252), .B(n233), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b9) );
  NOR2X1 U4582 ( .A(n179), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b0) );
  NOR2X1 U4583 ( .A(n200), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b0) );
  NOR2X1 U4584 ( .A(n242), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b0) );
  NOR2X1 U4585 ( .A(n270), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b0) );
  NOR2X1 U4586 ( .A(n199), .B(n4487), 
        .Y(input_p2_times_b2_mul_componentxUMxa15_and_b1) );
  NOR2X1 U4587 ( .A(n241), .B(n4593), 
        .Y(output_p2_times_a2_mul_componentxUMxa15_and_b1) );
  NOR2X1 U4588 ( .A(n194), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b6) );
  NOR2X1 U4589 ( .A(n236), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b6) );
  NOR2X1 U4590 ( .A(n179), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b0) );
  NOR2X1 U4591 ( .A(n200), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b0) );
  NOR2X1 U4592 ( .A(n242), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b0) );
  NOR2X1 U4593 ( .A(n270), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b0) );
  NOR2X1 U4594 ( .A(n172), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b7) );
  NOR2X1 U4595 ( .A(n193), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b7) );
  NOR2X1 U4596 ( .A(n235), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b7) );
  NOR2X1 U4597 ( .A(n263), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b7) );
  NOR2X1 U4598 ( .A(n170), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b9) );
  NOR2X1 U4599 ( .A(n261), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b9) );
  NOR2X1 U4600 ( .A(n171), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b8) );
  NOR2X1 U4601 ( .A(n262), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b8) );
  NOR2X1 U4602 ( .A(n191), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b9) );
  NOR2X1 U4603 ( .A(n233), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b9) );
  NOR2X1 U4604 ( .A(n192), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b8) );
  NOR2X1 U4605 ( .A(n234), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b8) );
  NOR2X1 U4606 ( .A(n178), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b1) );
  NOR2X1 U4607 ( .A(n199), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b1) );
  NOR2X1 U4608 ( .A(n241), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b1) );
  NOR2X1 U4609 ( .A(n269), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b1) );
  NOR2X1 U4610 ( .A(n171), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b8) );
  NOR2X1 U4611 ( .A(n192), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b8) );
  NOR2X1 U4612 ( .A(n234), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b8) );
  NOR2X1 U4613 ( .A(n262), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b8) );
  NOR2X1 U4614 ( .A(n180), .B(n173), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b6) );
  NOR2X1 U4615 ( .A(n201), .B(n194), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b6) );
  NOR2X1 U4616 ( .A(n243), .B(n236), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b6) );
  NOR2X1 U4617 ( .A(n271), .B(n264), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b6) );
  NOR2X1 U4618 ( .A(n180), .B(n172), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b7) );
  NOR2X1 U4619 ( .A(n201), .B(n193), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b7) );
  NOR2X1 U4620 ( .A(n243), .B(n235), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b7) );
  NOR2X1 U4621 ( .A(n271), .B(n263), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b7) );
  NOR2X1 U4622 ( .A(n175), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b4) );
  NOR2X1 U4623 ( .A(n196), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b4) );
  NOR2X1 U4624 ( .A(n238), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b4) );
  NOR2X1 U4625 ( .A(n266), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b4) );
  NOR2X1 U4626 ( .A(n195), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b5) );
  NOR2X1 U4627 ( .A(n237), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b5) );
  NOR2X1 U4628 ( .A(n174), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b5) );
  NOR2X1 U4629 ( .A(n195), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b5) );
  NOR2X1 U4630 ( .A(n237), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b5) );
  NOR2X1 U4631 ( .A(n265), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b5) );
  NOR2X1 U4632 ( .A(n173), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b6) );
  NOR2X1 U4633 ( .A(n194), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b6) );
  NOR2X1 U4634 ( .A(n236), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b6) );
  NOR2X1 U4635 ( .A(n264), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b6) );
  NOR2X1 U4636 ( .A(n173), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b6) );
  NOR2X1 U4637 ( .A(n194), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b6) );
  NOR2X1 U4638 ( .A(n236), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b6) );
  NOR2X1 U4639 ( .A(n264), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b6) );
  NOR2X1 U4640 ( .A(n173), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b6) );
  NOR2X1 U4641 ( .A(n194), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b6) );
  NOR2X1 U4642 ( .A(n236), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b6) );
  NOR2X1 U4643 ( .A(n264), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b6) );
  NOR2X1 U4644 ( .A(n172), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b7) );
  NOR2X1 U4645 ( .A(n263), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b7) );
  NOR2X1 U4646 ( .A(n170), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b9) );
  NOR2X1 U4647 ( .A(n261), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b9) );
  NOR2X1 U4648 ( .A(n171), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b8) );
  NOR2X1 U4649 ( .A(n262), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b8) );
  NOR2X1 U4650 ( .A(n193), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b7) );
  NOR2X1 U4651 ( .A(n235), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b7) );
  NOR2X1 U4652 ( .A(n191), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b9) );
  NOR2X1 U4653 ( .A(n233), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b9) );
  NOR2X1 U4654 ( .A(n192), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b8) );
  NOR2X1 U4655 ( .A(n234), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b8) );
  NOR2X1 U4656 ( .A(n172), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b7) );
  NOR2X1 U4657 ( .A(n193), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b7) );
  NOR2X1 U4658 ( .A(n235), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b7) );
  NOR2X1 U4659 ( .A(n263), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b7) );
  NOR2X1 U4660 ( .A(n171), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b8) );
  NOR2X1 U4661 ( .A(n192), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b8) );
  NOR2X1 U4662 ( .A(n234), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b8) );
  NOR2X1 U4663 ( .A(n262), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b8) );
  NOR2X1 U4664 ( .A(n170), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b9) );
  NOR2X1 U4665 ( .A(n261), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b9) );
  NOR2X1 U4666 ( .A(n191), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b9) );
  NOR2X1 U4667 ( .A(n233), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b9) );
  NOR2X1 U4668 ( .A(n175), .B(n4436), 
        .Y(input_p1_times_b1_mul_componentxUMxa13_and_b4) );
  NOR2X1 U4669 ( .A(n266), .B(input_times_b0_mul_componentxn85), 
        .Y(input_times_b0_mul_componentxUMxa13_and_b4) );
  NOR2X1 U4670 ( .A(n196), .B(n4489), 
        .Y(input_p2_times_b2_mul_componentxUMxa13_and_b4) );
  NOR2X1 U4671 ( .A(n238), .B(n4595), 
        .Y(output_p2_times_a2_mul_componentxUMxa13_and_b4) );
  NOR2X1 U4672 ( .A(n179), .B(n4433), 
        .Y(input_p1_times_b1_mul_componentxUMxa16_and_b0) );
  NOR2X1 U4673 ( .A(n270), .B(input_times_b0_mul_componentxn82), 
        .Y(input_times_b0_mul_componentxUMxa16_and_b0) );
  NOR2X1 U4674 ( .A(n200), .B(n4486), 
        .Y(input_p2_times_b2_mul_componentxUMxa16_and_b0) );
  NOR2X1 U4675 ( .A(n242), .B(n4592), 
        .Y(output_p2_times_a2_mul_componentxUMxa16_and_b0) );
  NOR2X1 U4676 ( .A(n179), .B(n10), 
        .Y(input_p1_times_b1_mul_componentxUMxa17_and_b0) );
  XOR2X1 U4677 ( .A(n3687), .B(input_previous_1[17]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[17]) );
  NOR2X1 U4678 ( .A(n200), .B(n11), 
        .Y(input_p2_times_b2_mul_componentxUMxa17_and_b0) );
  XOR2X1 U4679 ( .A(n3735), .B(input_previous_2[17]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[17]) );
  NOR2X1 U4680 ( .A(n242), .B(n12), 
        .Y(output_p2_times_a2_mul_componentxUMxa17_and_b0) );
  XOR2X1 U4681 ( .A(n3831), .B(output_previous_2[17]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[17]) );
  NOR2X1 U4682 ( .A(n270), .B(n13), 
        .Y(input_times_b0_mul_componentxUMxa17_and_b0) );
  XOR2X1 U4683 ( .A(n3639), .B(input_previous_0[17]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[17]) );
  XOR2X1 U4684 ( .A(input_p1_times_b1_mul_componentxUMxa15_and_b2), 
        .B(input_p1_times_b1_mul_componentxUMxa16_and_b1), .Y(n2718) );
  NOR2X1 U4685 ( .A(n177), .B(n4434), 
        .Y(input_p1_times_b1_mul_componentxUMxa15_and_b2) );
  NOR2X1 U4686 ( .A(n178), .B(n4433), 
        .Y(input_p1_times_b1_mul_componentxUMxa16_and_b1) );
  XOR2X1 U4687 ( .A(input_p1_times_b1_mul_componentxUMxa14_and_b3), .B(n2717), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127715984_127849024_127850928)
         );
  NOR2X1 U4688 ( .A(n176), .B(n4435), 
        .Y(input_p1_times_b1_mul_componentxUMxa14_and_b3) );
  XOR2X1 U4689 ( .A(input_p1_times_b1_mul_componentxUMxa12_and_b5), 
        .B(input_p1_times_b1_mul_componentxUMxa13_and_b4), .Y(n2717) );
  NOR2X1 U4690 ( .A(n174), .B(n4437), 
        .Y(input_p1_times_b1_mul_componentxUMxa12_and_b5) );
  XOR2X1 U4691 ( .A(input_p2_times_b2_mul_componentxUMxa15_and_b2), 
        .B(input_p2_times_b2_mul_componentxUMxa16_and_b1), .Y(n2952) );
  NOR2X1 U4692 ( .A(n198), .B(n4487), 
        .Y(input_p2_times_b2_mul_componentxUMxa15_and_b2) );
  NOR2X1 U4693 ( .A(n199), .B(n4486), 
        .Y(input_p2_times_b2_mul_componentxUMxa16_and_b1) );
  XOR2X1 U4694 ( .A(input_p2_times_b2_mul_componentxUMxa14_and_b3), .B(n2951), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127715984_127849024_127850928)
         );
  NOR2X1 U4695 ( .A(n197), .B(n4488), 
        .Y(input_p2_times_b2_mul_componentxUMxa14_and_b3) );
  XOR2X1 U4696 ( .A(input_p2_times_b2_mul_componentxUMxa12_and_b5), 
        .B(input_p2_times_b2_mul_componentxUMxa13_and_b4), .Y(n2951) );
  NOR2X1 U4697 ( .A(n195), .B(n4490), 
        .Y(input_p2_times_b2_mul_componentxUMxa12_and_b5) );
  XOR2X1 U4698 ( .A(output_p2_times_a2_mul_componentxUMxa15_and_b2), 
        .B(output_p2_times_a2_mul_componentxUMxa16_and_b1), .Y(n3420) );
  NOR2X1 U4699 ( .A(n240), .B(n4593), 
        .Y(output_p2_times_a2_mul_componentxUMxa15_and_b2) );
  NOR2X1 U4700 ( .A(n241), .B(n4592), 
        .Y(output_p2_times_a2_mul_componentxUMxa16_and_b1) );
  XOR2X1 U4701 ( .A(output_p2_times_a2_mul_componentxUMxa14_and_b3), .B(n3419), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127715984_127849024_127850928)
         );
  NOR2X1 U4702 ( .A(n239), .B(n4594), 
        .Y(output_p2_times_a2_mul_componentxUMxa14_and_b3) );
  XOR2X1 U4703 ( .A(output_p2_times_a2_mul_componentxUMxa12_and_b5), 
        .B(output_p2_times_a2_mul_componentxUMxa13_and_b4), .Y(n3419) );
  NOR2X1 U4704 ( .A(n237), .B(n4596), 
        .Y(output_p2_times_a2_mul_componentxUMxa12_and_b5) );
  XOR2X1 U4705 ( .A(input_times_b0_mul_componentxUMxa15_and_b2), 
        .B(input_times_b0_mul_componentxUMxa16_and_b1), .Y(n2484) );
  NOR2X1 U4706 ( .A(n268), .B(input_times_b0_mul_componentxn83), 
        .Y(input_times_b0_mul_componentxUMxa15_and_b2) );
  NOR2X1 U4707 ( .A(n269), .B(input_times_b0_mul_componentxn82), 
        .Y(input_times_b0_mul_componentxUMxa16_and_b1) );
  XOR2X1 U4708 ( .A(input_times_b0_mul_componentxUMxa14_and_b3), .B(n2483), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127715984_127849024_127850928)
         );
  NOR2X1 U4709 ( .A(n267), .B(input_times_b0_mul_componentxn84), 
        .Y(input_times_b0_mul_componentxUMxa14_and_b3) );
  XOR2X1 U4710 ( .A(input_times_b0_mul_componentxUMxa12_and_b5), 
        .B(input_times_b0_mul_componentxUMxa13_and_b4), .Y(n2483) );
  NOR2X1 U4711 ( .A(n265), .B(input_times_b0_mul_componentxn86), 
        .Y(input_times_b0_mul_componentxUMxa12_and_b5) );
  NOR2X1 U4712 ( .A(n4421), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b11) );
  NOR2X1 U4713 ( .A(n4474), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b11) );
  NOR2X1 U4714 ( .A(n4580), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b11) );
  NOR2X1 U4715 ( .A(input_times_b0_mul_componentxn70), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b11) );
  NOR2X1 U4716 ( .A(n4420), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b12) );
  NOR2X1 U4717 ( .A(n4473), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b12) );
  NOR2X1 U4718 ( .A(n4579), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b12) );
  NOR2X1 U4719 ( .A(input_times_b0_mul_componentxn69), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b12) );
  NOR2X1 U4720 ( .A(input_times_b0_mul_componentxn68), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b13) );
  NOR2X1 U4721 ( .A(n4419), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b13) );
  NOR2X1 U4722 ( .A(n4472), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b13) );
  NOR2X1 U4723 ( .A(n4578), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b13) );
  NOR2X1 U4724 ( .A(input_times_b0_mul_componentxn67), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b14) );
  NOR2X1 U4725 ( .A(n4418), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b14) );
  NOR2X1 U4726 ( .A(n4471), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b14) );
  NOR2X1 U4727 ( .A(n4577), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b14) );
  NOR2X1 U4728 ( .A(n4417), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b15) );
  NOR2X1 U4729 ( .A(n4470), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b15) );
  NOR2X1 U4730 ( .A(n4576), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b15) );
  NOR2X1 U4731 ( .A(input_times_b0_mul_componentxn66), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b15) );
  NOR2X1 U4732 ( .A(n192), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b8) );
  NOR2X1 U4733 ( .A(n234), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b8) );
  NOR2X1 U4734 ( .A(n170), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b9) );
  NOR2X1 U4735 ( .A(n191), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b9) );
  NOR2X1 U4736 ( .A(n233), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b9) );
  NOR2X1 U4737 ( .A(n261), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b9) );
  NOR2X1 U4738 ( .A(n4422), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b10) );
  NOR2X1 U4739 ( .A(n4475), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b10) );
  NOR2X1 U4740 ( .A(n4581), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b10) );
  NOR2X1 U4741 ( .A(input_times_b0_mul_componentxn71), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b10) );
  NOR2X1 U4742 ( .A(n4422), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b10) );
  NOR2X1 U4743 ( .A(n4475), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b10) );
  NOR2X1 U4744 ( .A(n4581), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b10) );
  NOR2X1 U4745 ( .A(input_times_b0_mul_componentxn71), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b10) );
  NOR2X1 U4746 ( .A(n4421), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b11) );
  NOR2X1 U4747 ( .A(n4474), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b11) );
  NOR2X1 U4748 ( .A(n4580), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b11) );
  NOR2X1 U4749 ( .A(input_times_b0_mul_componentxn70), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b11) );
  NOR2X1 U4750 ( .A(n4420), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b12) );
  NOR2X1 U4751 ( .A(n4473), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b12) );
  NOR2X1 U4752 ( .A(n4579), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b12) );
  NOR2X1 U4753 ( .A(input_times_b0_mul_componentxn69), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b12) );
  NOR2X1 U4754 ( .A(input_times_b0_mul_componentxn68), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b13) );
  NOR2X1 U4755 ( .A(n4420), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b12) );
  NOR2X1 U4756 ( .A(n4473), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b12) );
  NOR2X1 U4757 ( .A(n4579), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b12) );
  NOR2X1 U4758 ( .A(input_times_b0_mul_componentxn69), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b12) );
  NOR2X1 U4759 ( .A(n4419), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b13) );
  NOR2X1 U4760 ( .A(n4472), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b13) );
  NOR2X1 U4761 ( .A(n4578), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b13) );
  NOR2X1 U4762 ( .A(input_times_b0_mul_componentxn68), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b13) );
  NOR2X1 U4763 ( .A(n4419), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b13) );
  NOR2X1 U4764 ( .A(n4472), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b13) );
  NOR2X1 U4765 ( .A(n4578), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b13) );
  NOR2X1 U4766 ( .A(n280), .B(input_times_b0_mul_componentxn67), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b14) );
  NOR2X1 U4767 ( .A(n189), .B(n4418), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b14) );
  NOR2X1 U4768 ( .A(n210), .B(n4471), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b14) );
  NOR2X1 U4769 ( .A(n252), .B(n4577), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b14) );
  NOR2X1 U4770 ( .A(n189), .B(n4417), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b15) );
  NOR2X1 U4771 ( .A(n210), .B(n4470), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b15) );
  NOR2X1 U4772 ( .A(n252), .B(n4576), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b15) );
  NOR2X1 U4773 ( .A(n280), .B(input_times_b0_mul_componentxn66), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b15) );
  NOR2X1 U4774 ( .A(n189), .B(n4416), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b16) );
  NOR2X1 U4775 ( .A(n210), .B(n4469), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b16) );
  NOR2X1 U4776 ( .A(n252), .B(n4575), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b16) );
  NOR2X1 U4777 ( .A(n280), .B(input_times_b0_mul_componentxn65), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b16) );
  NOR2X1 U4778 ( .A(n170), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b9) );
  NOR2X1 U4779 ( .A(n261), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b9) );
  NOR2X1 U4780 ( .A(n191), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b9) );
  NOR2X1 U4781 ( .A(n233), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b9) );
  NOR2X1 U4782 ( .A(n172), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b7) );
  NOR2X1 U4783 ( .A(n193), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b7) );
  NOR2X1 U4784 ( .A(n235), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b7) );
  NOR2X1 U4785 ( .A(n263), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b7) );
  NOR2X1 U4786 ( .A(n171), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b8) );
  NOR2X1 U4787 ( .A(n192), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b8) );
  NOR2X1 U4788 ( .A(n234), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b8) );
  NOR2X1 U4789 ( .A(n262), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b8) );
  NOR2X1 U4790 ( .A(n189), .B(n178), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b1) );
  NOR2X1 U4791 ( .A(n280), .B(n269), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b1) );
  NOR2X1 U4792 ( .A(n210), .B(n199), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b1) );
  NOR2X1 U4793 ( .A(n252), .B(n241), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b1) );
  NOR2X1 U4794 ( .A(n179), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b0) );
  NOR2X1 U4795 ( .A(n200), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b0) );
  NOR2X1 U4796 ( .A(n242), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b0) );
  NOR2X1 U4797 ( .A(n270), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b0) );
  NOR2X1 U4798 ( .A(n173), .B(n4438), 
        .Y(input_p1_times_b1_mul_componentxUMxa11_and_b6) );
  NOR2X1 U4799 ( .A(n264), .B(input_times_b0_mul_componentxn87), 
        .Y(input_times_b0_mul_componentxUMxa11_and_b6) );
  NOR2X1 U4800 ( .A(n194), .B(n4491), 
        .Y(input_p2_times_b2_mul_componentxUMxa11_and_b6) );
  NOR2X1 U4801 ( .A(n236), .B(n4597), 
        .Y(output_p2_times_a2_mul_componentxUMxa11_and_b6) );
  XOR2X1 U4802 ( .A(input_p1_times_b1_mul_componentxUMxa9_and_b8), 
        .B(input_p1_times_b1_mul_componentxUMxa10_and_b7), .Y(n2716) );
  NOR2X1 U4803 ( .A(n180), .B(n171), 
        .Y(input_p1_times_b1_mul_componentxUMxa9_and_b8) );
  NOR2X1 U4804 ( .A(n172), .B(n4439), 
        .Y(input_p1_times_b1_mul_componentxUMxa10_and_b7) );
  XOR2X1 U4805 ( .A(input_p2_times_b2_mul_componentxUMxa9_and_b8), 
        .B(input_p2_times_b2_mul_componentxUMxa10_and_b7), .Y(n2950) );
  NOR2X1 U4806 ( .A(n201), .B(n192), 
        .Y(input_p2_times_b2_mul_componentxUMxa9_and_b8) );
  NOR2X1 U4807 ( .A(n193), .B(n4492), 
        .Y(input_p2_times_b2_mul_componentxUMxa10_and_b7) );
  XOR2X1 U4808 ( .A(output_p2_times_a2_mul_componentxUMxa9_and_b8), 
        .B(output_p2_times_a2_mul_componentxUMxa10_and_b7), .Y(n3418) );
  NOR2X1 U4809 ( .A(n243), .B(n234), 
        .Y(output_p2_times_a2_mul_componentxUMxa9_and_b8) );
  NOR2X1 U4810 ( .A(n235), .B(n4598), 
        .Y(output_p2_times_a2_mul_componentxUMxa10_and_b7) );
  XOR2X1 U4811 ( .A(input_times_b0_mul_componentxUMxa9_and_b8), 
        .B(input_times_b0_mul_componentxUMxa10_and_b7), .Y(n2482) );
  NOR2X1 U4812 ( .A(n271), .B(n262), 
        .Y(input_times_b0_mul_componentxUMxa9_and_b8) );
  NOR2X1 U4813 ( .A(n263), .B(input_times_b0_mul_componentxn88), 
        .Y(input_times_b0_mul_componentxUMxa10_and_b7) );
  XOR2X1 U4814 ( .A(input_p1_times_b1_mul_componentxUMxa6_and_b11), 
        .B(input_p1_times_b1_mul_componentxUMxa7_and_b10), .Y(n2715) );
  NOR2X1 U4815 ( .A(n4421), .B(n183), 
        .Y(input_p1_times_b1_mul_componentxUMxa6_and_b11) );
  NOR2X1 U4816 ( .A(n4422), .B(n182), 
        .Y(input_p1_times_b1_mul_componentxUMxa7_and_b10) );
  XOR2X1 U4817 ( .A(input_p2_times_b2_mul_componentxUMxa6_and_b11), 
        .B(input_p2_times_b2_mul_componentxUMxa7_and_b10), .Y(n2949) );
  NOR2X1 U4818 ( .A(n4474), .B(n204), 
        .Y(input_p2_times_b2_mul_componentxUMxa6_and_b11) );
  NOR2X1 U4819 ( .A(n4475), .B(n203), 
        .Y(input_p2_times_b2_mul_componentxUMxa7_and_b10) );
  XOR2X1 U4820 ( .A(output_p2_times_a2_mul_componentxUMxa6_and_b11), 
        .B(output_p2_times_a2_mul_componentxUMxa7_and_b10), .Y(n3417) );
  NOR2X1 U4821 ( .A(n4580), .B(n246), 
        .Y(output_p2_times_a2_mul_componentxUMxa6_and_b11) );
  NOR2X1 U4822 ( .A(n4581), .B(n245), 
        .Y(output_p2_times_a2_mul_componentxUMxa7_and_b10) );
  XOR2X1 U4823 ( .A(input_times_b0_mul_componentxUMxa6_and_b11), 
        .B(input_times_b0_mul_componentxUMxa7_and_b10), .Y(n2481) );
  NOR2X1 U4824 ( .A(input_times_b0_mul_componentxn70), .B(n274), 
        .Y(input_times_b0_mul_componentxUMxa6_and_b11) );
  NOR2X1 U4825 ( .A(input_times_b0_mul_componentxn71), .B(n273), 
        .Y(input_times_b0_mul_componentxUMxa7_and_b10) );
  NOR2X1 U4826 ( .A(n189), .B(n179), 
        .Y(input_p1_times_b1_mul_componentxUMxfirst_vector[0]) );
  NOR2X1 U4827 ( .A(n210), .B(n200), 
        .Y(input_p2_times_b2_mul_componentxUMxfirst_vector[0]) );
  NOR2X1 U4828 ( .A(n252), .B(n242), 
        .Y(output_p2_times_a2_mul_componentxUMxfirst_vector[0]) );
  NOR2X1 U4829 ( .A(n280), .B(n270), 
        .Y(input_times_b0_mul_componentxUMxfirst_vector[0]) );
  NOR2X1 U4830 ( .A(input_times_b0_mul_componentxn67), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b14) );
  NOR2X1 U4831 ( .A(n4418), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b14) );
  NOR2X1 U4832 ( .A(n4471), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b14) );
  NOR2X1 U4833 ( .A(n4577), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b14) );
  NOR2X1 U4834 ( .A(input_times_b0_mul_componentxn68), .B(n276), 
        .Y(input_times_b0_mul_componentxUMxa4_and_b13) );
  NOR2X1 U4835 ( .A(n4419), .B(n185), 
        .Y(input_p1_times_b1_mul_componentxUMxa4_and_b13) );
  NOR2X1 U4836 ( .A(n4472), .B(n206), 
        .Y(input_p2_times_b2_mul_componentxUMxa4_and_b13) );
  NOR2X1 U4837 ( .A(n4578), .B(n248), 
        .Y(output_p2_times_a2_mul_componentxUMxa4_and_b13) );
  NOR2X1 U4838 ( .A(n4417), .B(n187), 
        .Y(input_p1_times_b1_mul_componentxUMxa2_and_b15) );
  NOR2X1 U4839 ( .A(n4470), .B(n208), 
        .Y(input_p2_times_b2_mul_componentxUMxa2_and_b15) );
  NOR2X1 U4840 ( .A(n4576), .B(n250), 
        .Y(output_p2_times_a2_mul_componentxUMxa2_and_b15) );
  NOR2X1 U4841 ( .A(input_times_b0_mul_componentxn66), .B(n278), 
        .Y(input_times_b0_mul_componentxUMxa2_and_b15) );
  NOR2X1 U4842 ( .A(n170), .B(n181), 
        .Y(input_p1_times_b1_mul_componentxUMxa8_and_b9) );
  NOR2X1 U4843 ( .A(n191), .B(n202), 
        .Y(input_p2_times_b2_mul_componentxUMxa8_and_b9) );
  NOR2X1 U4844 ( .A(n233), .B(n244), 
        .Y(output_p2_times_a2_mul_componentxUMxa8_and_b9) );
  NOR2X1 U4845 ( .A(n261), .B(n272), 
        .Y(input_times_b0_mul_componentxUMxa8_and_b9) );
  XOR2X1 U4846 ( .A(input_p1_times_b1_mul_componentxUMxa0_and_b17), 
        .B(input_p1_times_b1_mul_componentxUMxa1_and_b16), .Y(n2713) );
  NOR2X1 U4847 ( .A(n189), .B(n21), 
        .Y(input_p1_times_b1_mul_componentxUMxa0_and_b17) );
  NOR2X1 U4848 ( .A(n4416), .B(n188), 
        .Y(input_p1_times_b1_mul_componentxUMxa1_and_b16) );
  XOR2X1 U4849 ( .A(input_p2_times_b2_mul_componentxUMxa0_and_b17), 
        .B(input_p2_times_b2_mul_componentxUMxa1_and_b16), .Y(n2947) );
  NOR2X1 U4850 ( .A(n210), .B(n22), 
        .Y(input_p2_times_b2_mul_componentxUMxa0_and_b17) );
  NOR2X1 U4851 ( .A(n4469), .B(n209), 
        .Y(input_p2_times_b2_mul_componentxUMxa1_and_b16) );
  XOR2X1 U4852 ( .A(output_p2_times_a2_mul_componentxUMxa0_and_b17), 
        .B(output_p2_times_a2_mul_componentxUMxa1_and_b16), .Y(n3415) );
  NOR2X1 U4853 ( .A(n252), .B(n23), 
        .Y(output_p2_times_a2_mul_componentxUMxa0_and_b17) );
  NOR2X1 U4854 ( .A(n4575), .B(n251), 
        .Y(output_p2_times_a2_mul_componentxUMxa1_and_b16) );
  XOR2X1 U4855 ( .A(input_times_b0_mul_componentxUMxa0_and_b17), 
        .B(input_times_b0_mul_componentxUMxa1_and_b16), .Y(n2479) );
  NOR2X1 U4856 ( .A(n280), .B(n24), 
        .Y(input_times_b0_mul_componentxUMxa0_and_b17) );
  NOR2X1 U4857 ( .A(input_times_b0_mul_componentxn65), .B(n279), 
        .Y(input_times_b0_mul_componentxUMxa1_and_b16) );
  XOR2X1 U4858 ( .A(input_p1_times_b1_mul_componentxUMxa5_and_b12), .B(n2714), 
        .Y(input_p1_times_b1_mul_componentxUMxsum_layer1_127674016_127675920_127731136)
         );
  NOR2X1 U4859 ( .A(n4420), .B(n184), 
        .Y(input_p1_times_b1_mul_componentxUMxa5_and_b12) );
  XOR2X1 U4860 ( .A(input_p1_times_b1_mul_componentxUMxa3_and_b14), 
        .B(input_p1_times_b1_mul_componentxUMxa4_and_b13), .Y(n2714) );
  NOR2X1 U4861 ( .A(n4418), .B(n186), 
        .Y(input_p1_times_b1_mul_componentxUMxa3_and_b14) );
  XOR2X1 U4862 ( .A(input_p2_times_b2_mul_componentxUMxa5_and_b12), .B(n2948), 
        .Y(input_p2_times_b2_mul_componentxUMxsum_layer1_127674016_127675920_127731136)
         );
  NOR2X1 U4863 ( .A(n4473), .B(n205), 
        .Y(input_p2_times_b2_mul_componentxUMxa5_and_b12) );
  XOR2X1 U4864 ( .A(input_p2_times_b2_mul_componentxUMxa3_and_b14), 
        .B(input_p2_times_b2_mul_componentxUMxa4_and_b13), .Y(n2948) );
  NOR2X1 U4865 ( .A(n4471), .B(n207), 
        .Y(input_p2_times_b2_mul_componentxUMxa3_and_b14) );
  XOR2X1 U4866 ( .A(output_p2_times_a2_mul_componentxUMxa5_and_b12), .B(n3416), 
        .Y(output_p2_times_a2_mul_componentxUMxsum_layer1_127674016_127675920_127731136)
         );
  NOR2X1 U4867 ( .A(n4579), .B(n247), 
        .Y(output_p2_times_a2_mul_componentxUMxa5_and_b12) );
  XOR2X1 U4868 ( .A(output_p2_times_a2_mul_componentxUMxa3_and_b14), 
        .B(output_p2_times_a2_mul_componentxUMxa4_and_b13), .Y(n3416) );
  NOR2X1 U4869 ( .A(n4577), .B(n249), 
        .Y(output_p2_times_a2_mul_componentxUMxa3_and_b14) );
  XOR2X1 U4870 ( .A(input_times_b0_mul_componentxUMxa5_and_b12), .B(n2480), 
        .Y(input_times_b0_mul_componentxUMxsum_layer1_127674016_127675920_127731136)
         );
  NOR2X1 U4871 ( .A(input_times_b0_mul_componentxn69), .B(n275), 
        .Y(input_times_b0_mul_componentxUMxa5_and_b12) );
  XOR2X1 U4872 ( .A(input_times_b0_mul_componentxUMxa3_and_b14), 
        .B(input_times_b0_mul_componentxUMxa4_and_b13), .Y(n2480) );
  NOR2X1 U4873 ( .A(input_times_b0_mul_componentxn67), .B(n277), 
        .Y(input_times_b0_mul_componentxUMxa3_and_b14) );
  OAI2BB2X1 U4874 ( .B0(n1174), .B1(n319), .A0N(input_previous_0[17]), 
        .A1N(n320), .Y(input_prev_0_registerxn20) );
  OR2X2 U4875 ( .A(n367), .B(change_input), .Y(n103) );
  INVX1 U4876 ( .A(n103), .Y(n1870) );
  OR2X2 U4877 ( .A(n367), .B(change_input), .Y(n104) );
  INVX1 U4878 ( .A(n104), .Y(n1980) );
  OR2X2 U4879 ( .A(n368), .B(change_input), .Y(n105) );
  INVX1 U4880 ( .A(n105), .Y(n2089) );
  OR2X2 U4881 ( .A(n368), .B(change_input), .Y(n106) );
  INVX1 U4882 ( .A(n106), .Y(n2199) );
  OR2X2 U4883 ( .A(n367), .B(change_input), .Y(n107) );
  INVX1 U4884 ( .A(n107), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn3) );
  INVX1 U4885 ( .A(change_input), .Y(n1260) );
  INVX1 U4886 ( .A(n4203), .Y(n374) );
  INVX1 U4887 ( .A(n4259), .Y(n376) );
  INVX1 U4888 ( .A(n4369), .Y(n378) );
  INVX1 U4889 ( .A(input_times_b0_div_componentxn24), .Y(n380) );
  AOI22X1 U4890 ( .A0(n335), .A1(n338), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_10_), .B1(n336), 
        .Y(n4422) );
  XOR2X1 U4891 ( .A(n3710), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_10_) );
  NAND2X1 U4892 ( .A(n3695), .B(n337), .Y(n3710) );
  AOI22X1 U4893 ( .A0(n326), .A1(n329), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_10_), .B1(n327), 
        .Y(n4475) );
  XOR2X1 U4894 ( .A(n3758), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_10_) );
  NAND2X1 U4895 ( .A(n3743), .B(n328), .Y(n3758) );
  AOI22X1 U4896 ( .A0(n362), .A1(n365), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_10_), .B1(n363), 
        .Y(n4528) );
  XOR2X1 U4897 ( .A(n3806), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_10_) );
  NAND2X1 U4898 ( .A(n3791), .B(n364), .Y(n3806) );
  AOI22X1 U4899 ( .A0(n353), .A1(n356), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_10_), .B1(n354), 
        .Y(n4581) );
  XOR2X1 U4900 ( .A(n3854), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_10_) );
  NAND2X1 U4901 ( .A(n3839), .B(n355), .Y(n3854) );
  AOI22X1 U4902 ( .A0(n344), .A1(n347), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_10_), .B1(n345), 
        .Y(input_times_b0_mul_componentxn71) );
  XOR2X1 U4903 ( .A(n3662), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_10_) );
  NAND2X1 U4904 ( .A(n3647), .B(n346), .Y(n3662) );
  AOI22X1 U4905 ( .A0(n362), .A1(n365), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_11_), .B1(n363), 
        .Y(n4527) );
  XOR2X1 U4906 ( .A(n3804), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_11_) );
  AOI22X1 U4907 ( .A0(n335), .A1(n338), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_11_), .B1(n336), 
        .Y(n4421) );
  XOR2X1 U4908 ( .A(n3708), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_11_) );
  AOI22X1 U4909 ( .A0(n326), .A1(n329), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_11_), .B1(n327), 
        .Y(n4474) );
  XOR2X1 U4910 ( .A(n3756), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_11_) );
  AOI22X1 U4911 ( .A0(n353), .A1(n356), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_11_), .B1(n354), 
        .Y(n4580) );
  XOR2X1 U4912 ( .A(n3852), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_11_) );
  AOI22X1 U4913 ( .A0(n344), .A1(n347), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_11_), .B1(n345), 
        .Y(input_times_b0_mul_componentxn70) );
  XOR2X1 U4914 ( .A(n3660), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_11_) );
  AOI22X1 U4915 ( .A0(n362), .A1(n364), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_12_), .B1(n363), 
        .Y(n4526) );
  XOR2X1 U4916 ( .A(n3805), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_12_) );
  OR2X2 U4917 ( .A(n3804), .B(n363), .Y(n3805) );
  AOI22X1 U4918 ( .A0(n335), .A1(n338), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_12_), .B1(n336), 
        .Y(n4420) );
  XOR2X1 U4919 ( .A(n3709), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_12_) );
  OR2X2 U4920 ( .A(n3708), .B(n336), .Y(n3709) );
  AOI22X1 U4921 ( .A0(n326), .A1(n329), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_12_), .B1(n327), 
        .Y(n4473) );
  XOR2X1 U4922 ( .A(n3757), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_12_) );
  OR2X2 U4923 ( .A(n3756), .B(n327), .Y(n3757) );
  AOI22X1 U4924 ( .A0(n353), .A1(n356), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_12_), .B1(n354), 
        .Y(n4579) );
  XOR2X1 U4925 ( .A(n3853), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_12_) );
  OR2X2 U4926 ( .A(n3852), .B(n354), .Y(n3853) );
  AOI22X1 U4927 ( .A0(n344), .A1(n347), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_12_), .B1(n345), 
        .Y(input_times_b0_mul_componentxn69) );
  XOR2X1 U4928 ( .A(n3661), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_12_) );
  OR2X2 U4929 ( .A(n3660), .B(n345), .Y(n3661) );
  AOI22X1 U4930 ( .A0(n341), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_9_), 
        .B1(\parameter_B0_div[7] ), .Y(input_times_b0_div_componentxn54) );
  XNOR2X1 U4931 ( .A(n3882), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_9_) );
  AOI22X1 U4932 ( .A0(n332), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_9_), 
        .B1(\parameter_B1_div[7] ), .Y(n4232) );
  XNOR2X1 U4933 ( .A(n3925), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_9_) );
  AOI22X1 U4934 ( .A0(n323), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_9_), 
        .B1(\parameter_B2_div[7] ), .Y(n4288) );
  XNOR2X1 U4935 ( .A(n3968), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_9_) );
  AOI22X1 U4936 ( .A0(n359), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_9_), 
        .B1(\parameter_A1_div[7] ), .Y(n4342) );
  XNOR2X1 U4937 ( .A(n4011), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_9_) );
  AOI22X1 U4938 ( .A0(n350), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_9_), 
        .B1(\parameter_A2_div[7] ), .Y(n4398) );
  XNOR2X1 U4939 ( .A(n4054), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_9_) );
  AOI22X1 U4940 ( .A0(n343), .A1(n348), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_13_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn68) );
  XOR2X1 U4941 ( .A(n3658), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_13_) );
  AOI22X1 U4942 ( .A0(n335), .A1(n339), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_13_), .B1(n336), 
        .Y(n4419) );
  XOR2X1 U4943 ( .A(n3706), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_13_) );
  AOI22X1 U4944 ( .A0(n326), .A1(n330), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_13_), .B1(n327), 
        .Y(n4472) );
  XOR2X1 U4945 ( .A(n3754), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_13_) );
  AOI22X1 U4946 ( .A0(n362), .A1(n364), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_13_), .B1(n363), 
        .Y(n4525) );
  XOR2X1 U4947 ( .A(n3802), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_13_) );
  AOI22X1 U4948 ( .A0(n353), .A1(n357), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_13_), .B1(n354), 
        .Y(n4578) );
  XOR2X1 U4949 ( .A(n3850), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_13_) );
  AOI22X1 U4950 ( .A0(n344), .A1(n348), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_14_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn67) );
  XOR2X1 U4951 ( .A(n3659), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_14_) );
  OR2X2 U4952 ( .A(n345), .B(n3658), .Y(n3659) );
  AOI22X1 U4953 ( .A0(n335), .A1(n339), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_14_), .B1(n336), 
        .Y(n4418) );
  XOR2X1 U4954 ( .A(n3707), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_14_) );
  OR2X2 U4955 ( .A(n336), .B(n3706), .Y(n3707) );
  AOI22X1 U4956 ( .A0(n326), .A1(n330), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_14_), .B1(n327), 
        .Y(n4471) );
  XOR2X1 U4957 ( .A(n3755), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_14_) );
  OR2X2 U4958 ( .A(n327), .B(n3754), .Y(n3755) );
  AOI22X1 U4959 ( .A0(n362), .A1(n366), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_14_), .B1(n363), 
        .Y(n4524) );
  XOR2X1 U4960 ( .A(n3803), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_14_) );
  OR2X2 U4961 ( .A(n363), .B(n3802), .Y(n3803) );
  AOI22X1 U4962 ( .A0(n353), .A1(n357), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_14_), .B1(n354), 
        .Y(n4577) );
  XOR2X1 U4963 ( .A(n3851), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_14_) );
  OR2X2 U4964 ( .A(n354), .B(n3850), .Y(n3851) );
  AOI22X1 U4965 ( .A0(n335), .A1(n337), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_15_), .B1(n335), 
        .Y(n4417) );
  XNOR2X1 U4966 ( .A(n3705), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_15_) );
  AOI22X1 U4967 ( .A0(n326), .A1(n328), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_15_), .B1(n326), 
        .Y(n4470) );
  XNOR2X1 U4968 ( .A(n3753), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_15_) );
  AOI22X1 U4969 ( .A0(n362), .A1(n364), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_15_), .B1(n362), 
        .Y(n4523) );
  XNOR2X1 U4970 ( .A(n3801), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_15_) );
  AOI22X1 U4971 ( .A0(n353), .A1(n355), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_15_), .B1(n353), 
        .Y(n4576) );
  XNOR2X1 U4972 ( .A(n3849), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_15_) );
  AOI22X1 U4973 ( .A0(n343), .A1(n346), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_15_), .B1(n345), 
        .Y(input_times_b0_mul_componentxn66) );
  XNOR2X1 U4974 ( .A(n3657), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_15_) );
  AOI22X1 U4975 ( .A0(n341), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_8_), .B1(n341), 
        .Y(input_times_b0_div_componentxn53) );
  XOR2X1 U4976 ( .A(n3883), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_8_) );
  OR2X2 U4977 ( .A(\parameter_B0_div[7] ), .B(n3884), .Y(n3883) );
  AOI22X1 U4978 ( .A0(n332), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_8_), .B1(n332), 
        .Y(n4231) );
  XOR2X1 U4979 ( .A(n3926), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_8_) );
  OR2X2 U4980 ( .A(\parameter_B1_div[7] ), .B(n3927), .Y(n3926) );
  AOI22X1 U4981 ( .A0(n323), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_8_), .B1(n323), 
        .Y(n4287) );
  XOR2X1 U4982 ( .A(n3969), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_8_) );
  OR2X2 U4983 ( .A(\parameter_B2_div[7] ), .B(n3970), .Y(n3969) );
  AOI22X1 U4984 ( .A0(n359), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_8_), .B1(n359), 
        .Y(n4341) );
  XOR2X1 U4985 ( .A(n4012), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_8_) );
  OR2X2 U4986 ( .A(\parameter_A1_div[7] ), .B(n4013), .Y(n4012) );
  AOI22X1 U4987 ( .A0(n350), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_8_), .B1(n350), 
        .Y(n4397) );
  XOR2X1 U4988 ( .A(n4055), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_8_) );
  OR2X2 U4989 ( .A(\parameter_A2_div[7] ), .B(n4056), .Y(n4055) );
  AOI22X1 U4990 ( .A0(n362), .A1(n364), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_16_), .B1(n362), 
        .Y(n4522) );
  XNOR2X1 U4991 ( .A(n3800), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_16_) );
  AOI22X1 U4992 ( .A0(n335), .A1(n337), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_16_), .B1(n335), 
        .Y(n4416) );
  XNOR2X1 U4993 ( .A(n3704), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_16_) );
  AOI22X1 U4994 ( .A0(n326), .A1(n328), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_16_), .B1(n326), 
        .Y(n4469) );
  XNOR2X1 U4995 ( .A(n3752), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_16_) );
  AOI22X1 U4996 ( .A0(n353), .A1(n355), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_16_), .B1(n353), 
        .Y(n4575) );
  XNOR2X1 U4997 ( .A(n3848), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_16_) );
  AOI22X1 U4998 ( .A0(n344), .A1(n346), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_16_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn65) );
  XNOR2X1 U4999 ( .A(n3656), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_16_) );
  AOI22X1 U5000 ( .A0(n341), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_7_), .B1(n341), 
        .Y(input_times_b0_div_componentxn52) );
  XOR2X1 U5001 ( .A(n3884), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_7_) );
  AOI22X1 U5002 ( .A0(n332), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_7_), .B1(n332), 
        .Y(n4230) );
  XOR2X1 U5003 ( .A(n3927), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_7_) );
  AOI22X1 U5004 ( .A0(n323), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_7_), .B1(n323), 
        .Y(n4286) );
  XOR2X1 U5005 ( .A(n3970), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_7_) );
  AOI22X1 U5006 ( .A0(n359), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_7_), .B1(n359), 
        .Y(n4340) );
  XOR2X1 U5007 ( .A(n4013), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_7_) );
  AOI22X1 U5008 ( .A0(n350), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_7_), .B1(n350), 
        .Y(n4396) );
  XOR2X1 U5009 ( .A(n4056), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_7_) );
  AOI22X1 U5010 ( .A0(n341), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_11_), .B1(n341), 
        .Y(input_times_b0_div_componentxn56) );
  XOR2X1 U5011 ( .A(n3895), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_11_) );
  AOI22X1 U5012 ( .A0(n332), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_11_), .B1(n332), 
        .Y(n4234) );
  XOR2X1 U5013 ( .A(n3938), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_11_) );
  AOI22X1 U5014 ( .A0(n323), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_11_), .B1(n323), 
        .Y(n4290) );
  XOR2X1 U5015 ( .A(n3981), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_11_) );
  AOI22X1 U5016 ( .A0(n359), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_11_), .B1(n359), 
        .Y(n4344) );
  XOR2X1 U5017 ( .A(n4024), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_11_) );
  AOI22X1 U5018 ( .A0(n350), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_11_), .B1(n350), 
        .Y(n4400) );
  XOR2X1 U5019 ( .A(n4067), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_11_) );
  AOI22X1 U5020 ( .A0(n341), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_13_), .B1(n341), 
        .Y(input_times_b0_div_componentxn58) );
  XOR2X1 U5021 ( .A(n3893), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_13_) );
  AOI22X1 U5022 ( .A0(n332), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_13_), .B1(n332), 
        .Y(n4236) );
  XOR2X1 U5023 ( .A(n3936), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_13_) );
  AOI22X1 U5024 ( .A0(n323), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_13_), .B1(n323), 
        .Y(n4292) );
  XOR2X1 U5025 ( .A(n3979), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_13_) );
  AOI22X1 U5026 ( .A0(n359), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_13_), .B1(n359), 
        .Y(n4346) );
  XOR2X1 U5027 ( .A(n4022), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_13_) );
  AOI22X1 U5028 ( .A0(n350), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_13_), .B1(n350), 
        .Y(n4402) );
  XOR2X1 U5029 ( .A(n4065), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_13_) );
  AOI22X1 U5030 ( .A0(n341), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_10_), 
        .B1(\parameter_B0_div[7] ), .Y(input_times_b0_div_componentxn55) );
  XOR2X1 U5031 ( .A(n3897), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_10_) );
  NAND2X1 U5032 ( .A(n3882), .B(n342), .Y(n3897) );
  AOI22X1 U5033 ( .A0(n332), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_10_), 
        .B1(\parameter_B1_div[7] ), .Y(n4233) );
  XOR2X1 U5034 ( .A(n3940), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_10_) );
  NAND2X1 U5035 ( .A(n3925), .B(n333), .Y(n3940) );
  AOI22X1 U5036 ( .A0(n323), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_10_), 
        .B1(\parameter_B2_div[7] ), .Y(n4289) );
  XOR2X1 U5037 ( .A(n3983), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_10_) );
  NAND2X1 U5038 ( .A(n3968), .B(n324), .Y(n3983) );
  AOI22X1 U5039 ( .A0(n359), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_10_), 
        .B1(\parameter_A1_div[7] ), .Y(n4343) );
  XOR2X1 U5040 ( .A(n4026), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_10_) );
  NAND2X1 U5041 ( .A(n4011), .B(n360), .Y(n4026) );
  AOI22X1 U5042 ( .A0(n350), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_10_), 
        .B1(\parameter_A2_div[7] ), .Y(n4399) );
  XOR2X1 U5043 ( .A(n4069), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_10_) );
  NAND2X1 U5044 ( .A(n4054), .B(n351), .Y(n4069) );
  AOI22X1 U5045 ( .A0(n341), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_12_), 
        .B1(\parameter_B0_div[7] ), .Y(input_times_b0_div_componentxn57) );
  XOR2X1 U5046 ( .A(n3896), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_12_) );
  OR2X2 U5047 ( .A(n3895), .B(\parameter_B0_div[7] ), .Y(n3896) );
  AOI22X1 U5048 ( .A0(n332), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_12_), 
        .B1(\parameter_B1_div[7] ), .Y(n4235) );
  XOR2X1 U5049 ( .A(n3939), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_12_) );
  OR2X2 U5050 ( .A(n3938), .B(\parameter_B1_div[7] ), .Y(n3939) );
  AOI22X1 U5051 ( .A0(n323), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_12_), 
        .B1(\parameter_B2_div[7] ), .Y(n4291) );
  XOR2X1 U5052 ( .A(n3982), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_12_) );
  OR2X2 U5053 ( .A(n3981), .B(\parameter_B2_div[7] ), .Y(n3982) );
  AOI22X1 U5054 ( .A0(n359), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_12_), 
        .B1(\parameter_A1_div[7] ), .Y(n4345) );
  XOR2X1 U5055 ( .A(n4025), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_12_) );
  OR2X2 U5056 ( .A(n4024), .B(\parameter_A1_div[7] ), .Y(n4025) );
  AOI22X1 U5057 ( .A0(n350), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_12_), 
        .B1(\parameter_A2_div[7] ), .Y(n4401) );
  XOR2X1 U5058 ( .A(n4068), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_12_) );
  OR2X2 U5059 ( .A(n4067), .B(\parameter_A2_div[7] ), .Y(n4068) );
  AOI22X1 U5060 ( .A0(n340), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_14_), 
        .B1(\parameter_B0_div[7] ), .Y(input_times_b0_div_componentxn59) );
  XOR2X1 U5061 ( .A(n3894), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_14_) );
  OR2X2 U5062 ( .A(\parameter_B0_div[7] ), .B(n3893), .Y(n3894) );
  AOI22X1 U5063 ( .A0(n331), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_14_), 
        .B1(\parameter_B1_div[7] ), .Y(n4237) );
  XOR2X1 U5064 ( .A(n3937), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_14_) );
  OR2X2 U5065 ( .A(\parameter_B1_div[7] ), .B(n3936), .Y(n3937) );
  AOI22X1 U5066 ( .A0(n322), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_14_), 
        .B1(\parameter_B2_div[7] ), .Y(n4293) );
  XOR2X1 U5067 ( .A(n3980), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_14_) );
  OR2X2 U5068 ( .A(\parameter_B2_div[7] ), .B(n3979), .Y(n3980) );
  AOI22X1 U5069 ( .A0(n358), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_14_), 
        .B1(\parameter_A1_div[7] ), .Y(n4347) );
  XOR2X1 U5070 ( .A(n4023), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_14_) );
  OR2X2 U5071 ( .A(\parameter_A1_div[7] ), .B(n4022), .Y(n4023) );
  AOI22X1 U5072 ( .A0(n349), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_14_), 
        .B1(\parameter_A2_div[7] ), .Y(n4403) );
  XOR2X1 U5073 ( .A(n4066), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_14_) );
  OR2X2 U5074 ( .A(\parameter_A2_div[7] ), .B(n4065), .Y(n4066) );
  AOI22X1 U5075 ( .A0(n340), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_15_), 
        .B1(\parameter_B0_div[7] ), .Y(input_times_b0_div_componentxn60) );
  XNOR2X1 U5076 ( .A(n3892), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_15_) );
  AOI22X1 U5077 ( .A0(n331), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_15_), 
        .B1(\parameter_B1_div[7] ), .Y(n4238) );
  XNOR2X1 U5078 ( .A(n3935), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_15_) );
  AOI22X1 U5079 ( .A0(n322), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_15_), 
        .B1(\parameter_B2_div[7] ), .Y(n4294) );
  XNOR2X1 U5080 ( .A(n3978), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_15_) );
  AOI22X1 U5081 ( .A0(n358), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_15_), 
        .B1(\parameter_A1_div[7] ), .Y(n4348) );
  XNOR2X1 U5082 ( .A(n4021), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_15_) );
  AOI22X1 U5083 ( .A0(n349), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_15_), 
        .B1(\parameter_A2_div[7] ), .Y(n4404) );
  XNOR2X1 U5084 ( .A(n4064), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_15_) );
  NOR2X1 U5085 ( .A(n336), .B(n3697), .Y(n3695) );
  NOR2X1 U5086 ( .A(n327), .B(n3745), .Y(n3743) );
  NOR2X1 U5087 ( .A(n363), .B(n3793), .Y(n3791) );
  NOR2X1 U5088 ( .A(n354), .B(n3841), .Y(n3839) );
  NOR2X1 U5089 ( .A(n345), .B(n3649), .Y(n3647) );
  NOR2X1 U5090 ( .A(\parameter_B0_div[7] ), .B(n3884), .Y(n3882) );
  NOR2X1 U5091 ( .A(\parameter_B1_div[7] ), .B(n3927), .Y(n3925) );
  NOR2X1 U5092 ( .A(\parameter_B2_div[7] ), .B(n3970), .Y(n3968) );
  NOR2X1 U5093 ( .A(\parameter_A1_div[7] ), .B(n4013), .Y(n4011) );
  NOR2X1 U5094 ( .A(\parameter_A2_div[7] ), .B(n4056), .Y(n4054) );
  NAND3BX1 U5095 ( .AN(n336), .B(n339), .C(n3695), .Y(n3708) );
  NAND3BX1 U5096 ( .AN(n327), .B(n330), .C(n3743), .Y(n3756) );
  NAND3BX1 U5097 ( .AN(n363), .B(n366), .C(n3791), .Y(n3804) );
  NAND3BX1 U5098 ( .AN(n354), .B(n357), .C(n3839), .Y(n3852) );
  NAND3BX1 U5099 ( .AN(n345), .B(n348), .C(n3647), .Y(n3660) );
  NAND3BX1 U5100 ( .AN(\parameter_B0_div[7] ), .B(n342), .C(n3882), .Y(n3895)
         );
  NAND3BX1 U5101 ( .AN(\parameter_B1_div[7] ), .B(n333), .C(n3925), .Y(n3938)
         );
  NAND3BX1 U5102 ( .AN(\parameter_B2_div[7] ), .B(n324), .C(n3968), .Y(n3981)
         );
  NAND3BX1 U5103 ( .AN(\parameter_A1_div[7] ), .B(n360), .C(n4011), .Y(n4024)
         );
  NAND3BX1 U5104 ( .AN(\parameter_A2_div[7] ), .B(n351), .C(n4054), .Y(n4067)
         );
  NOR2BX1 U5105 ( .AN(n3705), .B(n336), .Y(n3704) );
  NOR2BX1 U5106 ( .AN(n3753), .B(n327), .Y(n3752) );
  NOR2BX1 U5107 ( .AN(n3801), .B(n363), .Y(n3800) );
  NOR2BX1 U5108 ( .AN(n3849), .B(n354), .Y(n3848) );
  NOR2BX1 U5109 ( .AN(n3657), .B(n345), .Y(n3656) );
  NOR2X1 U5110 ( .A(n336), .B(n3706), .Y(n3705) );
  NOR2X1 U5111 ( .A(n327), .B(n3754), .Y(n3753) );
  NOR2X1 U5112 ( .A(n363), .B(n3802), .Y(n3801) );
  NOR2X1 U5113 ( .A(n354), .B(n3850), .Y(n3849) );
  NOR2X1 U5114 ( .A(n345), .B(n3658), .Y(n3657) );
  NOR2BX1 U5115 ( .AN(input_times_b0_div_componentxinput_B_inverted_17_), 
        .B(n342), .Y(input_times_b0_div_componentxunsigned_B_17) );
  XOR2X1 U5116 ( .A(n3890), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_17_) );
  NAND2BX1 U5117 ( .AN(\parameter_B0_div[7] ), .B(n3891), .Y(n3890) );
  NOR2BX1 U5118 ( .AN(input_p1_times_b1_div_componentxinput_B_inverted_17_), 
        .B(n333), .Y(input_p1_times_b1_div_componentxunsigned_B_17) );
  XOR2X1 U5119 ( .A(n3933), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_17_) );
  NAND2BX1 U5120 ( .AN(\parameter_B1_div[7] ), .B(n3934), .Y(n3933) );
  NOR2BX1 U5121 ( .AN(input_p2_times_b2_div_componentxinput_B_inverted_17_), 
        .B(n324), .Y(input_p2_times_b2_div_componentxunsigned_B_17) );
  XOR2X1 U5122 ( .A(n3976), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_17_) );
  NAND2BX1 U5123 ( .AN(\parameter_B2_div[7] ), .B(n3977), .Y(n3976) );
  NOR2BX1 U5124 ( .AN(output_p1_times_a1_div_componentxinput_B_inverted_17_), 
        .B(n360), .Y(output_p1_times_a1_div_componentxunsigned_B_17) );
  XOR2X1 U5125 ( .A(n4019), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_17_) );
  NAND2BX1 U5126 ( .AN(\parameter_A1_div[7] ), .B(n4020), .Y(n4019) );
  NOR2BX1 U5127 ( .AN(output_p2_times_a2_div_componentxinput_B_inverted_17_), 
        .B(n351), .Y(output_p2_times_a2_div_componentxunsigned_B_17) );
  XOR2X1 U5128 ( .A(n4062), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_17_) );
  NAND2BX1 U5129 ( .AN(\parameter_A2_div[7] ), .B(n4063), .Y(n4062) );
  OR2X2 U5130 ( .A(n3708), .B(n336), .Y(n3706) );
  OR2X2 U5131 ( .A(n3756), .B(n327), .Y(n3754) );
  OR2X2 U5132 ( .A(n3804), .B(n363), .Y(n3802) );
  OR2X2 U5133 ( .A(n3852), .B(n354), .Y(n3850) );
  OR2X2 U5134 ( .A(n3660), .B(n345), .Y(n3658) );
  XOR2X1 U5135 ( .A(n847), .B(n846), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[1]) );
  XOR2X1 U5136 ( .A(n1006), .B(n1005), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[1])
         );
  XOR2X1 U5137 ( .A(n1165), .B(n1164), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[1])
         );
  XOR2X1 U5138 ( .A(n529), .B(n528), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[1])
         );
  XOR2X1 U5139 ( .A(n688), .B(n687), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[1])
         );
  XNOR2X1 U5140 ( .A(n848), 
        .B(input_times_b0_div_componentxUDxinverter_for_substractionxn9), 
        .Y(input_times_b0_div_componentxUDxsub_ready_negative_divisor[2]) );
  NOR2X1 U5141 ( .A(n846), .B(n847), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn9) );
  XNOR2X1 U5142 ( .A(n1007), .B(n1765), 
        .Y(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[2])
         );
  NOR2X1 U5143 ( .A(n1005), .B(n1006), .Y(n1765) );
  XNOR2X1 U5144 ( .A(n1166), .B(n1774), 
        .Y(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[2])
         );
  NOR2X1 U5145 ( .A(n1164), .B(n1165), .Y(n1774) );
  XNOR2X1 U5146 ( .A(n530), .B(n1783), 
        .Y(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[2])
         );
  NOR2X1 U5147 ( .A(n528), .B(n529), .Y(n1783) );
  XNOR2X1 U5148 ( .A(n689), .B(n1792), 
        .Y(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[2])
         );
  NOR2X1 U5149 ( .A(n687), .B(n688), .Y(n1792) );
  INVX1 U5150 ( .A(n339), .Y(n335) );
  INVX1 U5151 ( .A(n330), .Y(n326) );
  INVX1 U5152 ( .A(n366), .Y(n362) );
  INVX1 U5153 ( .A(n357), .Y(n353) );
  INVX1 U5154 ( .A(n348), .Y(n344) );
  OR3XL U5155 ( .A(n847), .B(n848), .C(n846), 
        .Y(input_times_b0_div_componentxUDxinverter_for_substractionxn8) );
  OR3XL U5156 ( .A(n1006), .B(n1007), .C(n1005), .Y(n1764) );
  OR3XL U5157 ( .A(n1165), .B(n1166), .C(n1164), .Y(n1773) );
  OR3XL U5158 ( .A(n529), .B(n530), .C(n528), .Y(n1782) );
  OR3XL U5159 ( .A(n688), .B(n689), .C(n687), .Y(n1791) );
  INVX1 U5160 ( .A(n342), .Y(n341) );
  INVX1 U5161 ( .A(n333), .Y(n332) );
  INVX1 U5162 ( .A(n324), .Y(n323) );
  INVX1 U5163 ( .A(n360), .Y(n359) );
  INVX1 U5164 ( .A(n351), .Y(n350) );
  INVX1 U5165 ( .A(n339), .Y(n334) );
  INVX1 U5166 ( .A(n330), .Y(n325) );
  INVX1 U5167 ( .A(n357), .Y(n352) );
  INVX1 U5168 ( .A(n366), .Y(n361) );
  INVX1 U5169 ( .A(input_times_b0_div_componentxn48), .Y(n849) );
  INVX1 U5170 ( .A(n4226), .Y(n1008) );
  INVX1 U5171 ( .A(n4282), .Y(n1167) );
  INVX1 U5172 ( .A(n4336), .Y(n531) );
  INVX1 U5173 ( .A(n4392), .Y(n690) );
  INVX1 U5174 ( .A(input_times_b0_div_componentxn50), .Y(n851) );
  INVX1 U5175 ( .A(n4228), .Y(n1010) );
  INVX1 U5176 ( .A(n4284), .Y(n1169) );
  INVX1 U5177 ( .A(n4338), .Y(n533) );
  INVX1 U5178 ( .A(n4394), .Y(n692) );
  INVX1 U5179 ( .A(input_times_b0_div_componentxn49), .Y(n850) );
  INVX1 U5180 ( .A(n4227), .Y(n1009) );
  INVX1 U5181 ( .A(n4283), .Y(n1168) );
  INVX1 U5182 ( .A(n4337), .Y(n532) );
  INVX1 U5183 ( .A(n4393), .Y(n691) );
  INVX1 U5184 ( .A(input_times_b0_div_componentxn51), .Y(n852) );
  INVX1 U5185 ( .A(n4229), .Y(n1011) );
  INVX1 U5186 ( .A(n4285), .Y(n1170) );
  INVX1 U5187 ( .A(n4339), .Y(n534) );
  INVX1 U5188 ( .A(n4395), .Y(n693) );
  INVX1 U5189 ( .A(input_times_b0_div_componentxn61), .Y(n843) );
  AOI22X1 U5190 ( .A0(n340), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_16_), .B1(n341), 
        .Y(input_times_b0_div_componentxn61) );
  XNOR2X1 U5191 ( .A(n3891), .B(n340), 
        .Y(input_times_b0_div_componentxinput_B_inverted_16_) );
  INVX1 U5192 ( .A(n4239), .Y(n1002) );
  AOI22X1 U5193 ( .A0(n331), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_16_), .B1(n332), 
        .Y(n4239) );
  XNOR2X1 U5194 ( .A(n3934), .B(n331), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_16_) );
  INVX1 U5195 ( .A(n4295), .Y(n1161) );
  AOI22X1 U5196 ( .A0(n322), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_16_), .B1(n323), 
        .Y(n4295) );
  XNOR2X1 U5197 ( .A(n3977), .B(n322), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_16_) );
  INVX1 U5198 ( .A(n4349), .Y(n525) );
  AOI22X1 U5199 ( .A0(n358), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_16_), .B1(n359), 
        .Y(n4349) );
  XNOR2X1 U5200 ( .A(n4020), .B(n358), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_16_) );
  INVX1 U5201 ( .A(n4405), .Y(n684) );
  AOI22X1 U5202 ( .A0(n349), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_16_), .B1(n350), 
        .Y(n4405) );
  XNOR2X1 U5203 ( .A(n4063), .B(n349), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_16_) );
  XOR2X1 U5204 ( .A(n3703), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_17_) );
  NAND2BX1 U5205 ( .AN(n336), .B(n3704), .Y(n3703) );
  XOR2X1 U5206 ( .A(n3751), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_17_) );
  NAND2BX1 U5207 ( .AN(n327), .B(n3752), .Y(n3751) );
  XOR2X1 U5208 ( .A(n3847), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_17_) );
  NAND2BX1 U5209 ( .AN(n354), .B(n3848), .Y(n3847) );
  XOR2X1 U5210 ( .A(n3655), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_17_) );
  NAND2BX1 U5211 ( .AN(n345), .B(n3656), .Y(n3655) );
  INVX1 U5212 ( .A(input_times_b0_div_componentxn47), .Y(n848) );
  INVX1 U5213 ( .A(n4225), .Y(n1007) );
  INVX1 U5214 ( .A(n4281), .Y(n1166) );
  INVX1 U5215 ( .A(n4335), .Y(n530) );
  INVX1 U5216 ( .A(n4391), .Y(n689) );
  BUFX3 U5217 ( .A(n4409), .Y(n172) );
  AOI22X1 U5218 ( .A0(n335), .A1(n337), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_7_), .B1(n335), 
        .Y(n4409) );
  XOR2X1 U5219 ( .A(n3697), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_7_) );
  BUFX3 U5220 ( .A(n4462), .Y(n193) );
  AOI22X1 U5221 ( .A0(n326), .A1(n328), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_7_), .B1(n326), 
        .Y(n4462) );
  XOR2X1 U5222 ( .A(n3745), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_7_) );
  BUFX3 U5223 ( .A(n4515), .Y(n214) );
  AOI22X1 U5224 ( .A0(n362), .A1(n364), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_7_), .B1(n362), 
        .Y(n4515) );
  XOR2X1 U5225 ( .A(n3793), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_7_) );
  BUFX3 U5226 ( .A(n4568), .Y(n235) );
  AOI22X1 U5227 ( .A0(n353), .A1(n355), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_7_), .B1(n353), 
        .Y(n4568) );
  XOR2X1 U5228 ( .A(n3841), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_7_) );
  BUFX3 U5229 ( .A(input_times_b0_mul_componentxn58), .Y(n263) );
  AOI22X1 U5230 ( .A0(n344), .A1(n346), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_7_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn58) );
  XOR2X1 U5231 ( .A(n3649), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_7_) );
  BUFX3 U5232 ( .A(n4408), .Y(n171) );
  AOI22X1 U5233 ( .A0(n334), .A1(n337), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_8_), .B1(n335), 
        .Y(n4408) );
  XOR2X1 U5234 ( .A(n3696), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_8_) );
  OR2X2 U5235 ( .A(n336), .B(n3697), .Y(n3696) );
  BUFX3 U5236 ( .A(n4461), .Y(n192) );
  AOI22X1 U5237 ( .A0(n325), .A1(n328), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_8_), .B1(n326), 
        .Y(n4461) );
  XOR2X1 U5238 ( .A(n3744), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_8_) );
  OR2X2 U5239 ( .A(n327), .B(n3745), .Y(n3744) );
  BUFX3 U5240 ( .A(n4567), .Y(n234) );
  AOI22X1 U5241 ( .A0(n352), .A1(n355), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_8_), .B1(n353), 
        .Y(n4567) );
  XOR2X1 U5242 ( .A(n3840), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_8_) );
  OR2X2 U5243 ( .A(n354), .B(n3841), .Y(n3840) );
  BUFX3 U5244 ( .A(input_times_b0_mul_componentxn57), .Y(n262) );
  AOI22X1 U5245 ( .A0(n344), .A1(n346), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_8_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn57) );
  XOR2X1 U5246 ( .A(n3648), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_8_) );
  OR2X2 U5247 ( .A(n345), .B(n3649), .Y(n3648) );
  BUFX3 U5248 ( .A(n4514), .Y(n213) );
  AOI22X1 U5249 ( .A0(n361), .A1(n365), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_8_), .B1(n362), 
        .Y(n4514) );
  XOR2X1 U5250 ( .A(n3792), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_8_) );
  OR2X2 U5251 ( .A(n363), .B(n3793), .Y(n3792) );
  BUFX3 U5252 ( .A(n4407), .Y(n170) );
  AOI22X1 U5253 ( .A0(n334), .A1(n337), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_9_), .B1(n335), 
        .Y(n4407) );
  XNOR2X1 U5254 ( .A(n3695), .B(n334), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_9_) );
  BUFX3 U5255 ( .A(n4460), .Y(n191) );
  AOI22X1 U5256 ( .A0(n325), .A1(n328), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_9_), .B1(n326), 
        .Y(n4460) );
  XNOR2X1 U5257 ( .A(n3743), .B(n325), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_9_) );
  BUFX3 U5258 ( .A(n4566), .Y(n233) );
  AOI22X1 U5259 ( .A0(n352), .A1(n355), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_9_), .B1(n353), 
        .Y(n4566) );
  XNOR2X1 U5260 ( .A(n3839), .B(n352), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_9_) );
  BUFX3 U5261 ( .A(input_times_b0_mul_componentxn56), .Y(n261) );
  AOI22X1 U5262 ( .A0(n344), .A1(n346), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_9_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn56) );
  XNOR2X1 U5263 ( .A(n3647), .B(n343), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_9_) );
  BUFX3 U5264 ( .A(n4513), .Y(n212) );
  AOI22X1 U5265 ( .A0(n361), .A1(n366), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_9_), .B1(n362), 
        .Y(n4513) );
  XNOR2X1 U5266 ( .A(n3791), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_9_) );
  XOR2X1 U5267 ( .A(n3799), .B(n361), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_17_) );
  NAND2BX1 U5268 ( .AN(n363), .B(n3800), .Y(n3799) );
  INVX1 U5269 ( .A(n283), .Y(n317) );
  INVX1 U5270 ( .A(n301), .Y(n316) );
  INVX1 U5271 ( .A(n307), .Y(n318) );
  INVX1 U5272 ( .A(n308), .Y(n315) );
  BUFX3 U5273 ( .A(output_p2_times_a2_div_componentxoutput_sign_gated), 
        .Y(n169) );
  BUFX3 U5274 ( .A(output_p1_times_a1_div_componentxoutput_sign_gated), 
        .Y(n168) );
  BUFX3 U5275 ( .A(input_p1_times_b1_div_componentxoutput_sign_gated), 
        .Y(n166) );
  BUFX3 U5276 ( .A(input_times_b0_div_componentxoutput_sign_gated), .Y(n260)
         );
  INVX1 U5277 ( .A(n4359), .Y(n1311) );
  AOI22X1 U5278 ( .A0(output_p2_times_a2_div_componentxunsigned_output_1), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[1]), 
        .B1(n169), .Y(n4359) );
  XOR2X1 U5279 ( .A(output_p2_times_a2_div_componentxunsigned_output_1), 
        .B(output_p2_times_a2_div_componentxunsigned_output_inverted[0]), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[1]) );
  INVX1 U5280 ( .A(n4193), .Y(n1370) );
  AOI22X1 U5281 ( .A0(input_p1_times_b1_div_componentxunsigned_output_1), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[1]), 
        .B1(n166), .Y(n4193) );
  XOR2X1 U5282 ( .A(input_p1_times_b1_div_componentxunsigned_output_1), 
        .B(input_p1_times_b1_div_componentxunsigned_output_inverted[0]), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[1]) );
  OAI2BB1X1 U5283 ( 
        .A0N(output_p1_times_a1_div_componentxUDxshifted_substraction_result_0), 
        .A1N(n371), .B0(n2088), .Y(n2108) );
  AOI22X1 U5284 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_16), 
        .A1(n2089), .B0(output_p1_times_a1_div_componentxunsigned_A_17), 
        .B1(n2090), .Y(n2088) );
  NOR2BX1 U5285 ( .AN(output_p1_times_a1_div_componentxinput_A_inverted[17]), 
        .B(n232), .Y(output_p1_times_a1_div_componentxunsigned_A_17) );
  XOR2X1 U5286 ( .A(n4005), .B(n111), 
        .Y(output_p1_times_a1_div_componentxinput_A_inverted[17]) );
  OAI2BB1X1 U5287 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_1), 
        .B0(n2106), .Y(n2124) );
  AOI22X1 U5288 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_0), 
        .A1(n2089), .B0(n382), .B1(n2090), .Y(n2106) );
  INVX1 U5289 ( .A(n4317), .Y(n382) );
  AOI22X1 U5290 ( .A0(n517), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[1]), .B1(n112), 
        .Y(n4317) );
  OAI2BB1X1 U5291 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_2), 
        .B0(n2105), .Y(n2123) );
  AOI22X1 U5292 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_1), 
        .A1(n2089), .B0(n383), .B1(n2090), .Y(n2105) );
  INVX1 U5293 ( .A(n4318), .Y(n383) );
  AOI22X1 U5294 ( .A0(n516), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[2]), .B1(n112), 
        .Y(n4318) );
  OAI2BB1X1 U5295 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_3), 
        .B0(n2104), .Y(n2122) );
  AOI22X1 U5296 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_2), 
        .A1(n2089), .B0(n384), .B1(n2090), .Y(n2104) );
  INVX1 U5297 ( .A(n4319), .Y(n384) );
  AOI22X1 U5298 ( .A0(n509), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[3]), .B1(n112), 
        .Y(n4319) );
  OAI2BB1X1 U5299 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_4), 
        .B0(n2103), .Y(n2121) );
  AOI22X1 U5300 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_3), 
        .A1(n2089), .B0(n385), .B1(n2090), .Y(n2103) );
  INVX1 U5301 ( .A(n4320), .Y(n385) );
  AOI22X1 U5302 ( .A0(n503), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[4]), .B1(n112), 
        .Y(n4320) );
  OAI2BB1X1 U5303 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_5), 
        .B0(n2102), .Y(n2120) );
  AOI22X1 U5304 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_4), 
        .A1(n2089), .B0(n386), .B1(n2090), .Y(n2102) );
  INVX1 U5305 ( .A(n4321), .Y(n386) );
  AOI22X1 U5306 ( .A0(n495), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[5]), .B1(n112), 
        .Y(n4321) );
  OAI2BB1X1 U5307 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_6), 
        .B0(n2101), .Y(n2119) );
  AOI22X1 U5308 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_5), 
        .A1(n2089), .B0(n387), .B1(n2090), .Y(n2101) );
  INVX1 U5309 ( .A(n4322), .Y(n387) );
  AOI22X1 U5310 ( .A0(n488), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[6]), .B1(n112), 
        .Y(n4322) );
  OAI2BB1X1 U5311 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_7), 
        .B0(n2100), .Y(n2118) );
  AOI22X1 U5312 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_6), 
        .A1(n2089), .B0(n388), .B1(n2090), .Y(n2100) );
  INVX1 U5313 ( .A(n4323), .Y(n388) );
  AOI22X1 U5314 ( .A0(n480), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[7]), .B1(n112), 
        .Y(n4323) );
  OAI2BB1X1 U5315 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_8), 
        .B0(n2099), .Y(n2117) );
  AOI22X1 U5316 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_7), 
        .A1(n2089), .B0(n389), .B1(n2090), .Y(n2099) );
  INVX1 U5317 ( .A(n4324), .Y(n389) );
  AOI22X1 U5318 ( .A0(n473), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[8]), .B1(n112), 
        .Y(n4324) );
  OAI2BB1X1 U5319 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_9), 
        .B0(n2098), .Y(n2116) );
  AOI22X1 U5320 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_8), 
        .A1(n2089), .B0(n390), .B1(n2090), .Y(n2098) );
  INVX1 U5321 ( .A(n4325), .Y(n390) );
  AOI22X1 U5322 ( .A0(n463), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[9]), .B1(n111), 
        .Y(n4325) );
  OAI2BB1X1 U5323 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_10), 
        .B0(n2097), .Y(n2115) );
  AOI22X1 U5324 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_9), 
        .A1(n2089), .B0(n391), .B1(n2090), .Y(n2097) );
  INVX1 U5325 ( .A(n4326), .Y(n391) );
  AOI22X1 U5326 ( .A0(n453), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[10]), .B1(n111), 
        .Y(n4326) );
  OAI2BB1X1 U5327 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_11), 
        .B0(n2096), .Y(n2114) );
  AOI22X1 U5328 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_10), 
        .A1(n2089), .B0(n392), .B1(n2090), .Y(n2096) );
  INVX1 U5329 ( .A(n4327), .Y(n392) );
  AOI22X1 U5330 ( .A0(n441), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[11]), .B1(n111), 
        .Y(n4327) );
  OAI2BB1X1 U5331 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_12), 
        .B0(n2095), .Y(n2113) );
  AOI22X1 U5332 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_11), 
        .A1(n2089), .B0(n393), .B1(n2090), .Y(n2095) );
  INVX1 U5333 ( .A(n4328), .Y(n393) );
  AOI22X1 U5334 ( .A0(n432), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[12]), .B1(n111), 
        .Y(n4328) );
  OAI2BB1X1 U5335 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_13), 
        .B0(n2094), .Y(n2112) );
  AOI22XL U5336 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_12), 
        .A1(n2089), .B0(n394), .B1(n2090), .Y(n2094) );
  INVX1 U5337 ( .A(n4329), .Y(n394) );
  AOI22X1 U5338 ( .A0(n423), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[13]), .B1(n111), 
        .Y(n4329) );
  OAI2BB1X1 U5339 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_14), 
        .B0(n2093), .Y(n2111) );
  AOI22XL U5340 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_13), 
        .A1(n2089), .B0(n395), .B1(n2090), .Y(n2093) );
  INVX1 U5341 ( .A(n4330), .Y(n395) );
  AOI22X1 U5342 ( .A0(n417), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[14]), .B1(n111), 
        .Y(n4330) );
  OAI2BB1X1 U5343 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_15), 
        .B0(n2092), .Y(n2110) );
  AOI22XL U5344 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_14), 
        .A1(n2089), .B0(n396), .B1(n2090), .Y(n2092) );
  INVX1 U5345 ( .A(n4331), .Y(n396) );
  AOI22X1 U5346 ( .A0(n408), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[15]), .B1(n111), 
        .Y(n4331) );
  OAI2BB1X1 U5347 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_16), 
        .B0(n2091), .Y(n2109) );
  AOI22XL U5348 ( 
        .A0(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_15), 
        .A1(n2089), .B0(n397), .B1(n2090), .Y(n2091) );
  INVX1 U5349 ( .A(n4332), .Y(n397) );
  AOI22X1 U5350 ( .A0(n401), .A1(n232), 
        .B0(output_p1_times_a1_div_componentxinput_A_inverted[16]), .B1(n111), 
        .Y(n4332) );
  INVX1 U5351 ( .A(n4305), .Y(n1331) );
  AOI22X1 U5352 ( .A0(output_p1_times_a1_div_componentxunsigned_output_1), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[1]), 
        .B1(n168), .Y(n4305) );
  XOR2X1 U5353 ( .A(output_p1_times_a1_div_componentxunsigned_output_1), 
        .B(output_p1_times_a1_div_componentxunsigned_output_inverted[0]), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[1]) );
  INVX1 U5354 ( .A(input_times_b0_div_componentxn12), .Y(n1227) );
  AOI22X1 U5355 ( .A0(input_times_b0_div_componentxunsigned_output_1), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[1]), 
        .B1(n260), .Y(input_times_b0_div_componentxn12) );
  XOR2X1 U5356 ( .A(input_times_b0_div_componentxunsigned_output_1), 
        .B(input_times_b0_div_componentxunsigned_output_inverted[0]), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[1]) );
  NOR3X1 U5357 ( .A(input_p1_times_b1_div_componentxunsigned_output_7), 
        .B(input_p1_times_b1_div_componentxunsigned_output_8), .C(n3943), 
        .Y(n3941) );
  NOR3X1 U5358 ( .A(input_times_b0_div_componentxunsigned_output_7), 
        .B(input_times_b0_div_componentxunsigned_output_8), .C(n3900), 
        .Y(n3898) );
  NOR3X1 U5359 ( .A(output_p2_times_a2_div_componentxunsigned_output_7), 
        .B(output_p2_times_a2_div_componentxunsigned_output_8), .C(n4072), 
        .Y(n4070) );
  NOR3X1 U5360 ( .A(output_p1_times_a1_div_componentxunsigned_output_7), 
        .B(output_p1_times_a1_div_componentxunsigned_output_8), .C(n4029), 
        .Y(n4027) );
  INVX1 U5361 ( .A(n4303), .Y(n1329) );
  AOI22X1 U5362 ( .A0(output_p1_times_a1_div_componentxunsigned_output_3), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[3]), 
        .B1(n168), .Y(n4303) );
  XOR2X1 U5363 ( .A(n4033), 
        .B(output_p1_times_a1_div_componentxunsigned_output_3), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[3]) );
  INVX1 U5364 ( .A(input_times_b0_div_componentxn10), .Y(n1223) );
  AOI22X1 U5365 ( .A0(input_times_b0_div_componentxunsigned_output_3), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[3]), 
        .B1(n260), .Y(input_times_b0_div_componentxn10) );
  XOR2X1 U5366 ( .A(n3904), .B(input_times_b0_div_componentxunsigned_output_3), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[3]) );
  INVX1 U5367 ( .A(n4301), .Y(n1327) );
  AOI22X1 U5368 ( .A0(output_p1_times_a1_div_componentxunsigned_output_5), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[5]), 
        .B1(n168), .Y(n4301) );
  XOR2X1 U5369 ( .A(n4031), 
        .B(output_p1_times_a1_div_componentxunsigned_output_5), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[5]) );
  INVX1 U5370 ( .A(input_times_b0_div_componentxn8), .Y(n1219) );
  AOI22X1 U5371 ( .A0(input_times_b0_div_componentxunsigned_output_5), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[5]), 
        .B1(n260), .Y(input_times_b0_div_componentxn8) );
  XOR2X1 U5372 ( .A(n3902), .B(input_times_b0_div_componentxunsigned_output_5), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[5]) );
  INVX1 U5373 ( .A(n4299), .Y(n1325) );
  AOI22X1 U5374 ( .A0(output_p1_times_a1_div_componentxunsigned_output_7), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[7]), 
        .B1(n168), .Y(n4299) );
  XOR2X1 U5375 ( .A(n4029), 
        .B(output_p1_times_a1_div_componentxunsigned_output_7), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[7]) );
  INVX1 U5376 ( .A(input_times_b0_div_componentxn6), .Y(n1215) );
  AOI22X1 U5377 ( .A0(input_times_b0_div_componentxunsigned_output_7), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[7]), 
        .B1(n260), .Y(input_times_b0_div_componentxn6) );
  XOR2X1 U5378 ( .A(n3900), .B(input_times_b0_div_componentxunsigned_output_7), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[7]) );
  INVX1 U5379 ( .A(n4201), .Y(n1378) );
  AOI22X1 U5380 ( .A0(input_p1_times_b1_div_componentxunsigned_output_10), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[10]), 
        .B1(n166), .Y(n4201) );
  XOR2X1 U5381 ( .A(n3956), 
        .B(input_p1_times_b1_div_componentxunsigned_output_10), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[10]) );
  NAND2X1 U5382 ( .A(n3941), .B(n1448), .Y(n3956) );
  INVX1 U5383 ( .A(input_times_b0_div_componentxn17), .Y(n1232) );
  AOI22X1 U5384 ( .A0(input_times_b0_div_componentxunsigned_output_13), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[13]), 
        .B1(n260), .Y(input_times_b0_div_componentxn17) );
  XOR2X1 U5385 ( .A(n3909), 
        .B(input_times_b0_div_componentxunsigned_output_13), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[13]) );
  NAND3BX1 U5386 ( .AN(input_p1_times_b1_div_componentxunsigned_output_10), 
        .B(n1448), .C(n3941), .Y(n3954) );
  NAND3BX1 U5387 ( .AN(input_times_b0_div_componentxunsigned_output_10), 
        .B(n1272), .C(n3898), .Y(n3911) );
  OR3XL U5388 ( .A(output_p2_times_a2_div_componentxunsigned_output_5), 
        .B(output_p2_times_a2_div_componentxunsigned_output_6), .C(n4074), 
        .Y(n4072) );
  OR3XL U5389 ( .A(output_p1_times_a1_div_componentxunsigned_output_5), 
        .B(output_p1_times_a1_div_componentxunsigned_output_6), .C(n4031), 
        .Y(n4029) );
  OR3XL U5390 ( .A(input_p1_times_b1_div_componentxunsigned_output_5), 
        .B(input_p1_times_b1_div_componentxunsigned_output_6), .C(n3945), 
        .Y(n3943) );
  OR3XL U5391 ( .A(input_times_b0_div_componentxunsigned_output_5), 
        .B(input_times_b0_div_componentxunsigned_output_6), .C(n3902), 
        .Y(n3900) );
  OR3XL U5392 ( .A(input_p1_times_b1_div_componentxunsigned_output_11), 
        .B(input_p1_times_b1_div_componentxunsigned_output_12), .C(n3954), 
        .Y(n3952) );
  OR3XL U5393 ( .A(input_times_b0_div_componentxunsigned_output_11), 
        .B(input_times_b0_div_componentxunsigned_output_12), .C(n3911), 
        .Y(n3909) );
  BUFX3 U5394 ( .A(input_p2_times_b2_div_componentxoutput_sign_gated), 
        .Y(n167) );
  OR3XL U5395 ( .A(output_p2_times_a2_div_componentxunsigned_output_1), 
        .B(output_p2_times_a2_div_componentxunsigned_output_2), 
        .C(output_p2_times_a2_div_componentxunsigned_output_inverted[0]), 
        .Y(n4076) );
  OR3XL U5396 ( .A(output_p1_times_a1_div_componentxunsigned_output_1), 
        .B(output_p1_times_a1_div_componentxunsigned_output_2), 
        .C(output_p1_times_a1_div_componentxunsigned_output_inverted[0]), 
        .Y(n4033) );
  OR3XL U5397 ( .A(input_p1_times_b1_div_componentxunsigned_output_1), 
        .B(input_p1_times_b1_div_componentxunsigned_output_2), 
        .C(input_p1_times_b1_div_componentxunsigned_output_inverted[0]), 
        .Y(n3947) );
  OR3XL U5398 ( .A(input_times_b0_div_componentxunsigned_output_1), 
        .B(input_times_b0_div_componentxunsigned_output_2), 
        .C(input_times_b0_div_componentxunsigned_output_inverted[0]), 
        .Y(n3904) );
  OR3XL U5399 ( .A(input_p2_times_b2_div_componentxunsigned_output_1), 
        .B(input_p2_times_b2_div_componentxunsigned_output_2), 
        .C(input_p2_times_b2_div_componentxunsigned_output_inverted[0]), 
        .Y(n3990) );
  OR3XL U5400 ( .A(output_p2_times_a2_div_componentxunsigned_output_3), 
        .B(output_p2_times_a2_div_componentxunsigned_output_4), .C(n4076), 
        .Y(n4074) );
  OR3XL U5401 ( .A(output_p1_times_a1_div_componentxunsigned_output_3), 
        .B(output_p1_times_a1_div_componentxunsigned_output_4), .C(n4033), 
        .Y(n4031) );
  OR3XL U5402 ( .A(input_p1_times_b1_div_componentxunsigned_output_3), 
        .B(input_p1_times_b1_div_componentxunsigned_output_4), .C(n3947), 
        .Y(n3945) );
  OR3XL U5403 ( .A(input_times_b0_div_componentxunsigned_output_3), 
        .B(input_times_b0_div_componentxunsigned_output_4), .C(n3904), 
        .Y(n3902) );
  INVX1 U5404 ( .A(input_times_b0_div_componentxn21), .Y(n1237) );
  AOI22X1 U5405 ( 
        .A0(input_times_b0_div_componentxunsigned_output_inverted[0]), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[0]), 
        .B1(n260), .Y(input_times_b0_div_componentxn21) );
  INVX1 U5406 ( .A(n4314), .Y(n1340) );
  AOI22X1 U5407 ( 
        .A0(output_p1_times_a1_div_componentxunsigned_output_inverted[0]), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[0]), 
        .B1(n168), .Y(n4314) );
  INVX1 U5408 ( .A(n4357), .Y(n1309) );
  AOI22X1 U5409 ( .A0(output_p2_times_a2_div_componentxunsigned_output_3), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[3]), 
        .B1(n169), .Y(n4357) );
  XOR2X1 U5410 ( .A(n4076), 
        .B(output_p2_times_a2_div_componentxunsigned_output_3), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[3]) );
  INVX1 U5411 ( .A(n4191), .Y(n1368) );
  AOI22X1 U5412 ( .A0(input_p1_times_b1_div_componentxunsigned_output_3), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[3]), 
        .B1(n166), .Y(n4191) );
  XOR2X1 U5413 ( .A(n3947), 
        .B(input_p1_times_b1_div_componentxunsigned_output_3), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[3]) );
  INVX1 U5414 ( .A(n4355), .Y(n1307) );
  AOI22X1 U5415 ( .A0(output_p2_times_a2_div_componentxunsigned_output_5), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[5]), 
        .B1(n169), .Y(n4355) );
  XOR2X1 U5416 ( .A(n4074), 
        .B(output_p2_times_a2_div_componentxunsigned_output_5), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[5]) );
  INVX1 U5417 ( .A(n4247), .Y(n1348) );
  AOI22X1 U5418 ( .A0(input_p2_times_b2_div_componentxunsigned_output_3), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[3]), 
        .B1(n167), .Y(n4247) );
  XOR2X1 U5419 ( .A(n3990), 
        .B(input_p2_times_b2_div_componentxunsigned_output_3), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[3]) );
  INVX1 U5420 ( .A(n4189), .Y(n1366) );
  AOI22X1 U5421 ( .A0(input_p1_times_b1_div_componentxunsigned_output_5), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[5]), 
        .B1(n166), .Y(n4189) );
  XOR2X1 U5422 ( .A(n3945), 
        .B(input_p1_times_b1_div_componentxunsigned_output_5), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[5]) );
  INVX1 U5423 ( .A(n4353), .Y(n1305) );
  AOI22X1 U5424 ( .A0(output_p2_times_a2_div_componentxunsigned_output_7), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[7]), 
        .B1(n169), .Y(n4353) );
  XOR2X1 U5425 ( .A(n4072), 
        .B(output_p2_times_a2_div_componentxunsigned_output_7), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[7]) );
  INVX1 U5426 ( .A(n4187), .Y(n1364) );
  AOI22X1 U5427 ( .A0(input_p1_times_b1_div_componentxunsigned_output_7), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[7]), 
        .B1(n166), .Y(n4187) );
  XOR2X1 U5428 ( .A(n3943), 
        .B(input_p1_times_b1_div_componentxunsigned_output_7), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[7]) );
  INVX1 U5429 ( .A(n4351), .Y(n1303) );
  AOI22X1 U5430 ( .A0(output_p2_times_a2_div_componentxunsigned_output_9), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[9]), 
        .B1(n169), .Y(n4351) );
  XNOR2X1 U5431 ( .A(n4070), 
        .B(output_p2_times_a2_div_componentxunsigned_output_9), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[9]) );
  INVX1 U5432 ( .A(n4185), .Y(n1362) );
  AOI22X1 U5433 ( .A0(input_p1_times_b1_div_componentxunsigned_output_9), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[9]), 
        .B1(n166), .Y(n4185) );
  XNOR2X1 U5434 ( .A(n3941), 
        .B(input_p1_times_b1_div_componentxunsigned_output_9), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[9]) );
  INVX1 U5435 ( .A(n4198), .Y(n1375) );
  AOI22X1 U5436 ( .A0(input_p1_times_b1_div_componentxunsigned_output_13), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[13]), 
        .B1(n166), .Y(n4198) );
  XOR2X1 U5437 ( .A(n3952), 
        .B(input_p1_times_b1_div_componentxunsigned_output_13), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[13]) );
  INVX1 U5438 ( .A(n4202), .Y(n1379) );
  AOI22X1 U5439 ( 
        .A0(input_p1_times_b1_div_componentxunsigned_output_inverted[0]), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[0]), 
        .B1(n166), .Y(n4202) );
  INVX1 U5440 ( .A(n4368), .Y(n1320) );
  AOI22X1 U5441 ( 
        .A0(output_p2_times_a2_div_componentxunsigned_output_inverted[0]), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[0]), 
        .B1(n169), .Y(n4368) );
  INVX1 U5442 ( .A(n4258), .Y(n1359) );
  AOI22X1 U5443 ( 
        .A0(input_p2_times_b2_div_componentxunsigned_output_inverted[0]), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[0]), 
        .B1(n167), .Y(n4258) );
  INVX1 U5444 ( .A(n4200), .Y(n1377) );
  AOI22X1 U5445 ( .A0(input_p1_times_b1_div_componentxunsigned_output_11), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[11]), 
        .B1(n166), .Y(n4200) );
  XOR2X1 U5446 ( .A(n3954), 
        .B(input_p1_times_b1_div_componentxunsigned_output_11), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[11]) );
  INVX1 U5447 ( .A(input_times_b0_div_componentxn19), .Y(n1234) );
  AOI22X1 U5448 ( .A0(input_times_b0_div_componentxunsigned_output_11), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[11]), 
        .B1(n260), .Y(input_times_b0_div_componentxn19) );
  XOR2X1 U5449 ( .A(n3911), 
        .B(input_times_b0_div_componentxunsigned_output_11), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[11]) );
  INVX1 U5450 ( .A(n4249), .Y(n1350) );
  AOI22X1 U5451 ( .A0(input_p2_times_b2_div_componentxunsigned_output_1), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[1]), 
        .B1(n167), .Y(n4249) );
  XOR2X1 U5452 ( .A(input_p2_times_b2_div_componentxunsigned_output_1), 
        .B(input_p2_times_b2_div_componentxunsigned_output_inverted[0]), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[1]) );
  INVX1 U5453 ( .A(n4297), .Y(n1323) );
  AOI22X1 U5454 ( .A0(output_p1_times_a1_div_componentxunsigned_output_9), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[9]), 
        .B1(n168), .Y(n4297) );
  XNOR2X1 U5455 ( .A(n4027), 
        .B(output_p1_times_a1_div_componentxunsigned_output_9), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[9]) );
  INVX1 U5456 ( .A(input_times_b0_div_componentxn3), .Y(n1211) );
  AOI22X1 U5457 ( .A0(input_times_b0_div_componentxunsigned_output_9), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[9]), 
        .B1(n260), .Y(input_times_b0_div_componentxn3) );
  XNOR2X1 U5458 ( .A(n3898), 
        .B(input_times_b0_div_componentxunsigned_output_9), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[9]) );
  INVX1 U5459 ( .A(n4358), .Y(n1310) );
  AOI22X1 U5460 ( .A0(output_p2_times_a2_div_componentxunsigned_output_2), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[2]), 
        .B1(n169), .Y(n4358) );
  XNOR2X1 U5461 ( .A(output_p2_times_a2_div_componentxunsigned_output_2), 
        .B(n4077), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[2]) );
  NOR2X1 U5462 ( 
        .A(output_p2_times_a2_div_componentxunsigned_output_inverted[0]), 
        .B(output_p2_times_a2_div_componentxunsigned_output_1), .Y(n4077) );
  INVX1 U5463 ( .A(n4192), .Y(n1369) );
  AOI22X1 U5464 ( .A0(input_p1_times_b1_div_componentxunsigned_output_2), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[2]), 
        .B1(n166), .Y(n4192) );
  XNOR2X1 U5465 ( .A(input_p1_times_b1_div_componentxunsigned_output_2), 
        .B(n3948), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[2]) );
  NOR2X1 U5466 ( 
        .A(input_p1_times_b1_div_componentxunsigned_output_inverted[0]), 
        .B(input_p1_times_b1_div_componentxunsigned_output_1), .Y(n3948) );
  INVX1 U5467 ( .A(n4356), .Y(n1308) );
  AOI22X1 U5468 ( .A0(output_p2_times_a2_div_componentxunsigned_output_4), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[4]), 
        .B1(n169), .Y(n4356) );
  XOR2X1 U5469 ( .A(n4075), 
        .B(output_p2_times_a2_div_componentxunsigned_output_4), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[4]) );
  OR2X2 U5470 ( .A(output_p2_times_a2_div_componentxunsigned_output_3), 
        .B(n4076), .Y(n4075) );
  INVX1 U5471 ( .A(n4248), .Y(n1349) );
  AOI22X1 U5472 ( .A0(input_p2_times_b2_div_componentxunsigned_output_2), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[2]), 
        .B1(n167), .Y(n4248) );
  XNOR2X1 U5473 ( .A(input_p2_times_b2_div_componentxunsigned_output_2), 
        .B(n3991), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[2]) );
  NOR2X1 U5474 ( 
        .A(input_p2_times_b2_div_componentxunsigned_output_inverted[0]), 
        .B(input_p2_times_b2_div_componentxunsigned_output_1), .Y(n3991) );
  INVX1 U5475 ( .A(n4190), .Y(n1367) );
  AOI22X1 U5476 ( .A0(input_p1_times_b1_div_componentxunsigned_output_4), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[4]), 
        .B1(n166), .Y(n4190) );
  XOR2X1 U5477 ( .A(n3946), 
        .B(input_p1_times_b1_div_componentxunsigned_output_4), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[4]) );
  OR2X2 U5478 ( .A(input_p1_times_b1_div_componentxunsigned_output_3), 
        .B(n3947), .Y(n3946) );
  INVX1 U5479 ( .A(n4354), .Y(n1306) );
  AOI22X1 U5480 ( .A0(output_p2_times_a2_div_componentxunsigned_output_6), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[6]), 
        .B1(n169), .Y(n4354) );
  XOR2X1 U5481 ( .A(n4073), 
        .B(output_p2_times_a2_div_componentxunsigned_output_6), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[6]) );
  OR2X2 U5482 ( .A(output_p2_times_a2_div_componentxunsigned_output_5), 
        .B(n4074), .Y(n4073) );
  INVX1 U5483 ( .A(n4188), .Y(n1365) );
  AOI22X1 U5484 ( .A0(input_p1_times_b1_div_componentxunsigned_output_6), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[6]), 
        .B1(n166), .Y(n4188) );
  XOR2X1 U5485 ( .A(n3944), 
        .B(input_p1_times_b1_div_componentxunsigned_output_6), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[6]) );
  OR2X2 U5486 ( .A(input_p1_times_b1_div_componentxunsigned_output_5), 
        .B(n3945), .Y(n3944) );
  INVX1 U5487 ( .A(n4352), .Y(n1304) );
  AOI22X1 U5488 ( .A0(output_p2_times_a2_div_componentxunsigned_output_8), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[8]), 
        .B1(n169), .Y(n4352) );
  XOR2X1 U5489 ( .A(n4071), 
        .B(output_p2_times_a2_div_componentxunsigned_output_8), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[8]) );
  OR2X2 U5490 ( .A(output_p2_times_a2_div_componentxunsigned_output_7), 
        .B(n4072), .Y(n4071) );
  INVX1 U5491 ( .A(n4186), .Y(n1363) );
  AOI22X1 U5492 ( .A0(input_p1_times_b1_div_componentxunsigned_output_8), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[8]), 
        .B1(n166), .Y(n4186) );
  XOR2X1 U5493 ( .A(n3942), 
        .B(input_p1_times_b1_div_componentxunsigned_output_8), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[8]) );
  OR2X2 U5494 ( .A(input_p1_times_b1_div_componentxunsigned_output_7), 
        .B(n3943), .Y(n3942) );
  INVX1 U5495 ( .A(n4199), .Y(n1376) );
  AOI22X1 U5496 ( .A0(input_p1_times_b1_div_componentxunsigned_output_12), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[12]), 
        .B1(n166), .Y(n4199) );
  XOR2X1 U5497 ( .A(n3955), 
        .B(input_p1_times_b1_div_componentxunsigned_output_12), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[12]) );
  OR2X2 U5498 ( .A(n3954), 
        .B(input_p1_times_b1_div_componentxunsigned_output_11), .Y(n3955) );
  INVX1 U5499 ( .A(n4197), .Y(n1374) );
  AOI22X1 U5500 ( .A0(input_p1_times_b1_div_componentxunsigned_output_14), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[14]), 
        .B1(n166), .Y(n4197) );
  XOR2X1 U5501 ( .A(n3953), 
        .B(input_p1_times_b1_div_componentxunsigned_output_14), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[14]) );
  OR2X2 U5502 ( .A(input_p1_times_b1_div_componentxunsigned_output_13), 
        .B(n3952), .Y(n3953) );
  OAI2BB1X1 U5503 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_0), 
        .B0(n2107), .Y(n2125) );
  NAND2XL U5504 ( .A(n381), .B(n2090), .Y(n2107) );
  INVX1 U5505 ( .A(n4316), .Y(n381) );
  AOI22X1 U5506 ( .A0(n518), .A1(n232), .B0(n518), .B1(n112), .Y(n4316) );
  INVX1 U5507 ( .A(n4304), .Y(n1330) );
  AOI22X1 U5508 ( .A0(output_p1_times_a1_div_componentxunsigned_output_2), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[2]), 
        .B1(n168), .Y(n4304) );
  XNOR2X1 U5509 ( .A(output_p1_times_a1_div_componentxunsigned_output_2), 
        .B(n4034), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[2]) );
  NOR2X1 U5510 ( 
        .A(output_p1_times_a1_div_componentxunsigned_output_inverted[0]), 
        .B(output_p1_times_a1_div_componentxunsigned_output_1), .Y(n4034) );
  INVX1 U5511 ( .A(input_times_b0_div_componentxn11), .Y(n1225) );
  AOI22X1 U5512 ( .A0(input_times_b0_div_componentxunsigned_output_2), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[2]), 
        .B1(n260), .Y(input_times_b0_div_componentxn11) );
  XNOR2X1 U5513 ( .A(input_times_b0_div_componentxunsigned_output_2), 
        .B(n3905), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[2]) );
  NOR2X1 U5514 ( .A(input_times_b0_div_componentxunsigned_output_inverted[0]), 
        .B(input_times_b0_div_componentxunsigned_output_1), .Y(n3905) );
  INVX1 U5515 ( .A(n4302), .Y(n1328) );
  AOI22X1 U5516 ( .A0(output_p1_times_a1_div_componentxunsigned_output_4), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[4]), 
        .B1(n168), .Y(n4302) );
  XOR2X1 U5517 ( .A(n4032), 
        .B(output_p1_times_a1_div_componentxunsigned_output_4), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[4]) );
  OR2X2 U5518 ( .A(output_p1_times_a1_div_componentxunsigned_output_3), 
        .B(n4033), .Y(n4032) );
  INVX1 U5519 ( .A(input_times_b0_div_componentxn9), .Y(n1221) );
  AOI22X1 U5520 ( .A0(input_times_b0_div_componentxunsigned_output_4), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[4]), 
        .B1(n260), .Y(input_times_b0_div_componentxn9) );
  XOR2X1 U5521 ( .A(n3903), .B(input_times_b0_div_componentxunsigned_output_4), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[4]) );
  OR2X2 U5522 ( .A(input_times_b0_div_componentxunsigned_output_3), .B(n3904), 
        .Y(n3903) );
  INVX1 U5523 ( .A(n4300), .Y(n1326) );
  AOI22X1 U5524 ( .A0(output_p1_times_a1_div_componentxunsigned_output_6), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[6]), 
        .B1(n168), .Y(n4300) );
  XOR2X1 U5525 ( .A(n4030), 
        .B(output_p1_times_a1_div_componentxunsigned_output_6), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[6]) );
  OR2X2 U5526 ( .A(output_p1_times_a1_div_componentxunsigned_output_5), 
        .B(n4031), .Y(n4030) );
  INVX1 U5527 ( .A(input_times_b0_div_componentxn7), .Y(n1217) );
  AOI22X1 U5528 ( .A0(input_times_b0_div_componentxunsigned_output_6), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[6]), 
        .B1(n260), .Y(input_times_b0_div_componentxn7) );
  XOR2X1 U5529 ( .A(n3901), .B(input_times_b0_div_componentxunsigned_output_6), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[6]) );
  OR2X2 U5530 ( .A(input_times_b0_div_componentxunsigned_output_5), .B(n3902), 
        .Y(n3901) );
  INVX1 U5531 ( .A(n4298), .Y(n1324) );
  AOI22X1 U5532 ( .A0(output_p1_times_a1_div_componentxunsigned_output_8), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[8]), 
        .B1(n168), .Y(n4298) );
  XOR2X1 U5533 ( .A(n4028), 
        .B(output_p1_times_a1_div_componentxunsigned_output_8), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[8]) );
  OR2X2 U5534 ( .A(output_p1_times_a1_div_componentxunsigned_output_7), 
        .B(n4029), .Y(n4028) );
  INVX1 U5535 ( .A(input_times_b0_div_componentxn5), .Y(n1213) );
  AOI22X1 U5536 ( .A0(input_times_b0_div_componentxunsigned_output_8), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[8]), 
        .B1(n260), .Y(input_times_b0_div_componentxn5) );
  XOR2X1 U5537 ( .A(n3899), .B(input_times_b0_div_componentxunsigned_output_8), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[8]) );
  OR2X2 U5538 ( .A(input_times_b0_div_componentxunsigned_output_7), .B(n3900), 
        .Y(n3899) );
  INVX1 U5539 ( .A(input_times_b0_div_componentxn20), .Y(n1235) );
  AOI22X1 U5540 ( .A0(input_times_b0_div_componentxunsigned_output_10), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[10]), 
        .B1(n260), .Y(input_times_b0_div_componentxn20) );
  XOR2X1 U5541 ( .A(n3913), 
        .B(input_times_b0_div_componentxunsigned_output_10), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[10]) );
  NAND2X1 U5542 ( .A(n3898), .B(n1272), .Y(n3913) );
  INVX1 U5543 ( .A(input_times_b0_div_componentxn18), .Y(n1233) );
  AOI22X1 U5544 ( .A0(input_times_b0_div_componentxunsigned_output_12), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[12]), 
        .B1(n260), .Y(input_times_b0_div_componentxn18) );
  XOR2X1 U5545 ( .A(n3912), 
        .B(input_times_b0_div_componentxunsigned_output_12), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[12]) );
  OR2X2 U5546 ( .A(n3911), .B(input_times_b0_div_componentxunsigned_output_11), 
        .Y(n3912) );
  OAI2BB2X1 U5547 ( .B0(n108), .B1(n147), .A0N(n4315), .A1N(n108), .Y(n4350)
         );
  AND2X2 U5548 ( .A(output_p1_times_a1_div_componentxoutput_ready_signal), 
        .B(en), .Y(n108) );
  NOR3X1 U5549 ( .A(input_p2_times_b2_div_componentxunsigned_output_7), 
        .B(input_p2_times_b2_div_componentxunsigned_output_8), .C(n3986), 
        .Y(n3984) );
  NOR3X1 U5550 ( .A(input_p1_times_b1_div_componentxunsigned_output_13), 
        .B(input_p1_times_b1_div_componentxunsigned_output_14), .C(n3952), 
        .Y(n3951) );
  NOR3X1 U5551 ( .A(input_times_b0_div_componentxunsigned_output_13), 
        .B(input_times_b0_div_componentxunsigned_output_14), .C(n3909), 
        .Y(n3908) );
  NOR3X1 U5552 ( .A(output_p2_times_a2_div_componentxunsigned_output_13), 
        .B(output_p2_times_a2_div_componentxunsigned_output_14), .C(n4081), 
        .Y(n4080) );
  NOR3X1 U5553 ( .A(output_p1_times_a1_div_componentxunsigned_output_13), 
        .B(output_p1_times_a1_div_componentxunsigned_output_14), .C(n4038), 
        .Y(n4037) );
  NOR3X1 U5554 ( .A(input_p2_times_b2_div_componentxunsigned_output_13), 
        .B(input_p2_times_b2_div_componentxunsigned_output_14), .C(n3995), 
        .Y(n3994) );
  INVX1 U5555 ( .A(n4367), .Y(n1319) );
  AOI22X1 U5556 ( .A0(output_p2_times_a2_div_componentxunsigned_output_10), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[10]), 
        .B1(n169), .Y(n4367) );
  XOR2X1 U5557 ( .A(n4085), 
        .B(output_p2_times_a2_div_componentxunsigned_output_10), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[10]) );
  NAND2X1 U5558 ( .A(n4070), .B(n1391), .Y(n4085) );
  INVX1 U5559 ( .A(n4257), .Y(n1358) );
  AOI22X1 U5560 ( .A0(input_p2_times_b2_div_componentxunsigned_output_10), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[10]), 
        .B1(n167), .Y(n4257) );
  XOR2X1 U5561 ( .A(n3999), 
        .B(input_p2_times_b2_div_componentxunsigned_output_10), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[10]) );
  NAND2X1 U5562 ( .A(n3984), .B(n1429), .Y(n3999) );
  INVX1 U5563 ( .A(n4310), .Y(n1336) );
  AOI22X1 U5564 ( .A0(output_p1_times_a1_div_componentxunsigned_output_13), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[13]), 
        .B1(n168), .Y(n4310) );
  XOR2X1 U5565 ( .A(n4038), 
        .B(output_p1_times_a1_div_componentxunsigned_output_13), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[13]) );
  AOI22X1 U5566 ( .A0(input_p1_times_b1_div_componentxunsigned_output_17), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[17]), 
        .B1(n166), .Y(n4194) );
  XOR2X1 U5567 ( .A(n3949), 
        .B(input_p1_times_b1_div_componentxunsigned_output_17), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[17]) );
  NAND2BX1 U5568 ( .AN(input_p1_times_b1_div_componentxunsigned_output_16), 
        .B(n3950), .Y(n3949) );
  NAND3BX1 U5569 ( .AN(output_p2_times_a2_div_componentxunsigned_output_10), 
        .B(n1391), .C(n4070), .Y(n4083) );
  NAND3BX1 U5570 ( .AN(output_p1_times_a1_div_componentxunsigned_output_10), 
        .B(n1410), .C(n4027), .Y(n4040) );
  NAND3BX1 U5571 ( .AN(input_p2_times_b2_div_componentxunsigned_output_10), 
        .B(n1429), .C(n3984), .Y(n3997) );
  NOR2BX1 U5572 ( .AN(n3951), 
        .B(input_p1_times_b1_div_componentxunsigned_output_15), .Y(n3950) );
  NOR2BX1 U5573 ( .AN(n3908), 
        .B(input_times_b0_div_componentxunsigned_output_15), .Y(n3907) );
  NOR2BX1 U5574 ( .AN(n4037), 
        .B(output_p1_times_a1_div_componentxunsigned_output_15), .Y(n4036) );
  NOR2BX1 U5575 ( .AN(n4080), 
        .B(output_p2_times_a2_div_componentxunsigned_output_15), .Y(n4079) );
  NOR2BX1 U5576 ( .AN(n3994), 
        .B(input_p2_times_b2_div_componentxunsigned_output_15), .Y(n3993) );
  OR3XL U5577 ( .A(input_p2_times_b2_div_componentxunsigned_output_5), 
        .B(input_p2_times_b2_div_componentxunsigned_output_6), .C(n3988), 
        .Y(n3986) );
  OR3XL U5578 ( .A(output_p2_times_a2_div_componentxunsigned_output_11), 
        .B(output_p2_times_a2_div_componentxunsigned_output_12), .C(n4083), 
        .Y(n4081) );
  OR3XL U5579 ( .A(output_p1_times_a1_div_componentxunsigned_output_11), 
        .B(output_p1_times_a1_div_componentxunsigned_output_12), .C(n4040), 
        .Y(n4038) );
  OR3XL U5580 ( .A(input_p2_times_b2_div_componentxunsigned_output_11), 
        .B(input_p2_times_b2_div_componentxunsigned_output_12), .C(n3997), 
        .Y(n3995) );
  OR3XL U5581 ( .A(input_p2_times_b2_div_componentxunsigned_output_3), 
        .B(input_p2_times_b2_div_componentxunsigned_output_4), .C(n3990), 
        .Y(n3988) );
  INVX1 U5582 ( .A(n4245), .Y(n1346) );
  AOI22X1 U5583 ( .A0(input_p2_times_b2_div_componentxunsigned_output_5), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[5]), 
        .B1(n167), .Y(n4245) );
  XOR2X1 U5584 ( .A(n3988), 
        .B(input_p2_times_b2_div_componentxunsigned_output_5), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[5]) );
  INVX1 U5585 ( .A(n4243), .Y(n1344) );
  AOI22X1 U5586 ( .A0(input_p2_times_b2_div_componentxunsigned_output_7), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[7]), 
        .B1(n167), .Y(n4243) );
  XOR2X1 U5587 ( .A(n3986), 
        .B(input_p2_times_b2_div_componentxunsigned_output_7), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[7]) );
  INVX1 U5588 ( .A(n4241), .Y(n1342) );
  AOI22X1 U5589 ( .A0(input_p2_times_b2_div_componentxunsigned_output_9), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[9]), 
        .B1(n167), .Y(n4241) );
  XNOR2X1 U5590 ( .A(n3984), 
        .B(input_p2_times_b2_div_componentxunsigned_output_9), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[9]) );
  INVX1 U5591 ( .A(n4364), .Y(n1316) );
  AOI22X1 U5592 ( .A0(output_p2_times_a2_div_componentxunsigned_output_13), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[13]), 
        .B1(n169), .Y(n4364) );
  XOR2X1 U5593 ( .A(n4081), 
        .B(output_p2_times_a2_div_componentxunsigned_output_13), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[13]) );
  INVX1 U5594 ( .A(n4254), .Y(n1355) );
  AOI22X1 U5595 ( .A0(input_p2_times_b2_div_componentxunsigned_output_13), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[13]), 
        .B1(n167), .Y(n4254) );
  XOR2X1 U5596 ( .A(n3995), 
        .B(input_p2_times_b2_div_componentxunsigned_output_13), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[13]) );
  INVX1 U5597 ( .A(n4196), .Y(n1373) );
  AOI22X1 U5598 ( .A0(input_p1_times_b1_div_componentxunsigned_output_15), 
        .A1(n151), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[15]), 
        .B1(n166), .Y(n4196) );
  XNOR2X1 U5599 ( .A(n3951), 
        .B(input_p1_times_b1_div_componentxunsigned_output_15), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[15]) );
  INVX1 U5600 ( .A(n4362), .Y(n1314) );
  AOI22X1 U5601 ( .A0(output_p2_times_a2_div_componentxunsigned_output_15), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[15]), 
        .B1(n169), .Y(n4362) );
  XNOR2X1 U5602 ( .A(n4080), 
        .B(output_p2_times_a2_div_componentxunsigned_output_15), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[15]) );
  INVX1 U5603 ( .A(n4252), .Y(n1353) );
  AOI22X1 U5604 ( .A0(input_p2_times_b2_div_componentxunsigned_output_15), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[15]), 
        .B1(n167), .Y(n4252) );
  XNOR2X1 U5605 ( .A(n3994), 
        .B(input_p2_times_b2_div_componentxunsigned_output_15), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[15]) );
  INVX1 U5606 ( .A(n4195), .Y(n1372) );
  AOI22X1 U5607 ( .A0(input_p1_times_b1_div_componentxunsigned_output_16), 
        .A1(n152), 
        .B0(input_p1_times_b1_div_componentxunsigned_output_inverted[16]), 
        .B1(n166), .Y(n4195) );
  XNOR2X1 U5608 ( .A(n3950), 
        .B(input_p1_times_b1_div_componentxunsigned_output_16), 
        .Y(input_p1_times_b1_div_componentxunsigned_output_inverted[16]) );
  INVX1 U5609 ( .A(n4361), .Y(n1313) );
  AOI22X1 U5610 ( .A0(output_p2_times_a2_div_componentxunsigned_output_16), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[16]), 
        .B1(n169), .Y(n4361) );
  XNOR2X1 U5611 ( .A(n4079), 
        .B(output_p2_times_a2_div_componentxunsigned_output_16), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[16]) );
  INVX1 U5612 ( .A(n4251), .Y(n1352) );
  AOI22X1 U5613 ( .A0(input_p2_times_b2_div_componentxunsigned_output_16), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[16]), 
        .B1(n167), .Y(n4251) );
  XNOR2X1 U5614 ( .A(n3993), 
        .B(input_p2_times_b2_div_componentxunsigned_output_16), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[16]) );
  INVX1 U5615 ( .A(n4366), .Y(n1318) );
  AOI22X1 U5616 ( .A0(output_p2_times_a2_div_componentxunsigned_output_11), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[11]), 
        .B1(n169), .Y(n4366) );
  XOR2X1 U5617 ( .A(n4083), 
        .B(output_p2_times_a2_div_componentxunsigned_output_11), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[11]) );
  INVX1 U5618 ( .A(n4312), .Y(n1338) );
  AOI22X1 U5619 ( .A0(output_p1_times_a1_div_componentxunsigned_output_11), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[11]), 
        .B1(n168), .Y(n4312) );
  XOR2X1 U5620 ( .A(n4040), 
        .B(output_p1_times_a1_div_componentxunsigned_output_11), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[11]) );
  INVX1 U5621 ( .A(n4256), .Y(n1357) );
  AOI22X1 U5622 ( .A0(input_p2_times_b2_div_componentxunsigned_output_11), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[11]), 
        .B1(n167), .Y(n4256) );
  XOR2X1 U5623 ( .A(n3997), 
        .B(input_p2_times_b2_div_componentxunsigned_output_11), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[11]) );
  INVX1 U5624 ( .A(input_times_b0_div_componentxn15), .Y(n1230) );
  AOI22X1 U5625 ( .A0(input_times_b0_div_componentxunsigned_output_15), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[15]), 
        .B1(n260), .Y(input_times_b0_div_componentxn15) );
  XNOR2X1 U5626 ( .A(n3908), 
        .B(input_times_b0_div_componentxunsigned_output_15), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[15]) );
  INVX1 U5627 ( .A(n4308), .Y(n1334) );
  AOI22X1 U5628 ( .A0(output_p1_times_a1_div_componentxunsigned_output_15), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[15]), 
        .B1(n168), .Y(n4308) );
  XNOR2X1 U5629 ( .A(n4037), 
        .B(output_p1_times_a1_div_componentxunsigned_output_15), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[15]) );
  INVX1 U5630 ( .A(n4246), .Y(n1347) );
  AOI22X1 U5631 ( .A0(input_p2_times_b2_div_componentxunsigned_output_4), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[4]), 
        .B1(n167), .Y(n4246) );
  XOR2X1 U5632 ( .A(n3989), 
        .B(input_p2_times_b2_div_componentxunsigned_output_4), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[4]) );
  OR2X2 U5633 ( .A(input_p2_times_b2_div_componentxunsigned_output_3), 
        .B(n3990), .Y(n3989) );
  INVX1 U5634 ( .A(n4244), .Y(n1345) );
  AOI22X1 U5635 ( .A0(input_p2_times_b2_div_componentxunsigned_output_6), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[6]), 
        .B1(n167), .Y(n4244) );
  XOR2X1 U5636 ( .A(n3987), 
        .B(input_p2_times_b2_div_componentxunsigned_output_6), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[6]) );
  OR2X2 U5637 ( .A(input_p2_times_b2_div_componentxunsigned_output_5), 
        .B(n3988), .Y(n3987) );
  INVX1 U5638 ( .A(n4242), .Y(n1343) );
  AOI22X1 U5639 ( .A0(input_p2_times_b2_div_componentxunsigned_output_8), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[8]), 
        .B1(n167), .Y(n4242) );
  XOR2X1 U5640 ( .A(n3985), 
        .B(input_p2_times_b2_div_componentxunsigned_output_8), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[8]) );
  OR2X2 U5641 ( .A(input_p2_times_b2_div_componentxunsigned_output_7), 
        .B(n3986), .Y(n3985) );
  INVX1 U5642 ( .A(n4365), .Y(n1317) );
  AOI22X1 U5643 ( .A0(output_p2_times_a2_div_componentxunsigned_output_12), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[12]), 
        .B1(n169), .Y(n4365) );
  XOR2X1 U5644 ( .A(n4084), 
        .B(output_p2_times_a2_div_componentxunsigned_output_12), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[12]) );
  OR2X2 U5645 ( .A(n4083), 
        .B(output_p2_times_a2_div_componentxunsigned_output_11), .Y(n4084) );
  INVX1 U5646 ( .A(n4255), .Y(n1356) );
  AOI22X1 U5647 ( .A0(input_p2_times_b2_div_componentxunsigned_output_12), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[12]), 
        .B1(n167), .Y(n4255) );
  XOR2X1 U5648 ( .A(n3998), 
        .B(input_p2_times_b2_div_componentxunsigned_output_12), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[12]) );
  OR2X2 U5649 ( .A(n3997), 
        .B(input_p2_times_b2_div_componentxunsigned_output_11), .Y(n3998) );
  INVX1 U5650 ( .A(n4363), .Y(n1315) );
  AOI22X1 U5651 ( .A0(output_p2_times_a2_div_componentxunsigned_output_14), 
        .A1(n146), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[14]), 
        .B1(n169), .Y(n4363) );
  XOR2X1 U5652 ( .A(n4082), 
        .B(output_p2_times_a2_div_componentxunsigned_output_14), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[14]) );
  OR2X2 U5653 ( .A(output_p2_times_a2_div_componentxunsigned_output_13), 
        .B(n4081), .Y(n4082) );
  INVX1 U5654 ( .A(n4253), .Y(n1354) );
  AOI22X1 U5655 ( .A0(input_p2_times_b2_div_componentxunsigned_output_14), 
        .A1(n150), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[14]), 
        .B1(n167), .Y(n4253) );
  XOR2X1 U5656 ( .A(n3996), 
        .B(input_p2_times_b2_div_componentxunsigned_output_14), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[14]) );
  OR2X2 U5657 ( .A(input_p2_times_b2_div_componentxunsigned_output_13), 
        .B(n3995), .Y(n3996) );
  INVX1 U5658 ( .A(input_times_b0_div_componentxn14), .Y(n1229) );
  AOI22X1 U5659 ( .A0(input_times_b0_div_componentxunsigned_output_16), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[16]), 
        .B1(n260), .Y(input_times_b0_div_componentxn14) );
  XNOR2X1 U5660 ( .A(n3907), 
        .B(input_times_b0_div_componentxunsigned_output_16), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[16]) );
  INVX1 U5661 ( .A(n4307), .Y(n1333) );
  AOI22X1 U5662 ( .A0(output_p1_times_a1_div_componentxunsigned_output_16), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[16]), 
        .B1(n168), .Y(n4307) );
  XNOR2X1 U5663 ( .A(n4036), 
        .B(output_p1_times_a1_div_componentxunsigned_output_16), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[16]) );
  INVX1 U5664 ( .A(n4313), .Y(n1339) );
  AOI22X1 U5665 ( .A0(output_p1_times_a1_div_componentxunsigned_output_10), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[10]), 
        .B1(n168), .Y(n4313) );
  XOR2X1 U5666 ( .A(n4042), 
        .B(output_p1_times_a1_div_componentxunsigned_output_10), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[10]) );
  NAND2X1 U5667 ( .A(n4027), .B(n1410), .Y(n4042) );
  INVX1 U5668 ( .A(n4311), .Y(n1337) );
  AOI22X1 U5669 ( .A0(output_p1_times_a1_div_componentxunsigned_output_12), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[12]), 
        .B1(n168), .Y(n4311) );
  XOR2X1 U5670 ( .A(n4041), 
        .B(output_p1_times_a1_div_componentxunsigned_output_12), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[12]) );
  OR2X2 U5671 ( .A(n4040), 
        .B(output_p1_times_a1_div_componentxunsigned_output_11), .Y(n4041) );
  INVX1 U5672 ( .A(input_times_b0_div_componentxn16), .Y(n1231) );
  AOI22X1 U5673 ( .A0(input_times_b0_div_componentxunsigned_output_14), 
        .A1(n136), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[14]), 
        .B1(n260), .Y(input_times_b0_div_componentxn16) );
  XOR2X1 U5674 ( .A(n3910), 
        .B(input_times_b0_div_componentxunsigned_output_14), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[14]) );
  OR2X2 U5675 ( .A(input_times_b0_div_componentxunsigned_output_13), .B(n3909), 
        .Y(n3910) );
  INVX1 U5676 ( .A(n4309), .Y(n1335) );
  AOI22X1 U5677 ( .A0(output_p1_times_a1_div_componentxunsigned_output_14), 
        .A1(n148), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[14]), 
        .B1(n168), .Y(n4309) );
  XOR2X1 U5678 ( .A(n4039), 
        .B(output_p1_times_a1_div_componentxunsigned_output_14), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[14]) );
  OR2X2 U5679 ( .A(output_p1_times_a1_div_componentxunsigned_output_13), 
        .B(n4038), .Y(n4039) );
  INVX1 U5680 ( .A(input_times_b0_div_componentxn13), .Y(n1228) );
  AOI22X1 U5681 ( .A0(input_times_b0_div_componentxunsigned_output_17), 
        .A1(n135), 
        .B0(input_times_b0_div_componentxunsigned_output_inverted[17]), 
        .B1(n260), .Y(input_times_b0_div_componentxn13) );
  XOR2X1 U5682 ( .A(n3906), 
        .B(input_times_b0_div_componentxunsigned_output_17), 
        .Y(input_times_b0_div_componentxunsigned_output_inverted[17]) );
  NAND2BX1 U5683 ( .AN(input_times_b0_div_componentxunsigned_output_16), 
        .B(n3907), .Y(n3906) );
  INVX1 U5684 ( .A(n4306), .Y(n1332) );
  AOI22X1 U5685 ( .A0(output_p1_times_a1_div_componentxunsigned_output_17), 
        .A1(n147), 
        .B0(output_p1_times_a1_div_componentxunsigned_output_inverted[17]), 
        .B1(n168), .Y(n4306) );
  XOR2X1 U5686 ( .A(n4035), 
        .B(output_p1_times_a1_div_componentxunsigned_output_17), 
        .Y(output_p1_times_a1_div_componentxunsigned_output_inverted[17]) );
  NAND2BX1 U5687 ( .AN(output_p1_times_a1_div_componentxunsigned_output_16), 
        .B(n4036), .Y(n4035) );
  INVX1 U5688 ( .A(n4360), .Y(n1312) );
  AOI22X1 U5689 ( .A0(output_p2_times_a2_div_componentxunsigned_output_17), 
        .A1(n145), 
        .B0(output_p2_times_a2_div_componentxunsigned_output_inverted[17]), 
        .B1(n169), .Y(n4360) );
  XOR2X1 U5690 ( .A(n4078), 
        .B(output_p2_times_a2_div_componentxunsigned_output_17), 
        .Y(output_p2_times_a2_div_componentxunsigned_output_inverted[17]) );
  NAND2BX1 U5691 ( .AN(output_p2_times_a2_div_componentxunsigned_output_16), 
        .B(n4079), .Y(n4078) );
  AOI22X1 U5692 ( .A0(input_p2_times_b2_div_componentxunsigned_output_17), 
        .A1(n149), 
        .B0(input_p2_times_b2_div_componentxunsigned_output_inverted[17]), 
        .B1(n167), .Y(n4250) );
  XOR2X1 U5693 ( .A(n3992), 
        .B(input_p2_times_b2_div_componentxunsigned_output_17), 
        .Y(input_p2_times_b2_div_componentxunsigned_output_inverted[17]) );
  NAND2BX1 U5694 ( .AN(input_p2_times_b2_div_componentxunsigned_output_16), 
        .B(n3993), .Y(n3992) );
  INVX1 U5695 ( .A(input_p1_times_b1_div_componentxunsigned_output_9), 
        .Y(n1448) );
  INVX1 U5696 ( .A(input_times_b0_div_componentxunsigned_output_9), .Y(n1272)
         );
  INVX1 U5697 ( .A(output_p2_times_a2_div_componentxunsigned_output_9), 
        .Y(n1391) );
  INVX1 U5698 ( .A(output_p1_times_a1_div_componentxunsigned_output_9), 
        .Y(n1410) );
  INVX1 U5699 ( .A(input_p2_times_b2_div_componentxunsigned_output_9), 
        .Y(n1429) );
  AOI22X1 U5700 ( .A0(input_previous_1[10]), .A1(n143), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[10]), 
        .B1(input_previous_1[17]), .Y(n4439) );
  XOR2X1 U5701 ( .A(n3694), .B(input_previous_1[10]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[10]) );
  NAND2X1 U5702 ( .A(n3679), .B(n1293), .Y(n3694) );
  AOI22X1 U5703 ( .A0(input_previous_2[10]), .A1(n141), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[10]), 
        .B1(input_previous_2[17]), .Y(n4492) );
  XOR2X1 U5704 ( .A(n3742), .B(input_previous_2[10]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[10]) );
  NAND2X1 U5705 ( .A(n3727), .B(n1283), .Y(n3742) );
  AOI22X1 U5706 ( .A0(output_previous_2[10]), .A1(n139), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[10]), 
        .B1(output_previous_2[17]), .Y(n4598) );
  XOR2X1 U5707 ( .A(n3838), .B(output_previous_2[10]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[10]) );
  NAND2X1 U5708 ( .A(n3823), .B(n1282), .Y(n3838) );
  AOI22X1 U5709 ( .A0(input_previous_0[10]), .A1(n131), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[10]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn88) );
  XOR2X1 U5710 ( .A(n3646), .B(input_previous_0[10]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[10]) );
  NAND2X1 U5711 ( .A(n3631), .B(n1191), .Y(n3646) );
  AOI22X1 U5712 ( .A0(input_previous_1[11]), .A1(n143), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[11]), 
        .B1(input_previous_1[17]), .Y(n4438) );
  XOR2X1 U5713 ( .A(n3692), .B(input_previous_1[11]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[11]) );
  AOI22X1 U5714 ( .A0(input_previous_0[11]), .A1(n131), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[11]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn87) );
  XOR2X1 U5715 ( .A(n3644), .B(input_previous_0[11]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[11]) );
  NOR3X1 U5716 ( .A(input_previous_1[7]), .B(input_previous_1[8]), .C(n3681), 
        .Y(n3679) );
  NOR3X1 U5717 ( .A(input_previous_0[7]), .B(input_previous_0[8]), .C(n3633), 
        .Y(n3631) );
  NOR3X1 U5718 ( .A(input_previous_2[7]), .B(input_previous_2[8]), .C(n3729), 
        .Y(n3727) );
  NOR3X1 U5719 ( .A(output_previous_2[7]), .B(output_previous_2[8]), .C(n3825), 
        .Y(n3823) );
  NAND3BX1 U5720 ( .AN(input_previous_1[10]), .B(n1293), .C(n3679), .Y(n3692)
         );
  NAND3BX1 U5721 ( .AN(input_previous_0[10]), .B(n1191), .C(n3631), .Y(n3644)
         );
  OR3XL U5722 ( .A(input_previous_1[5]), .B(input_previous_1[6]), .C(n3683), 
        .Y(n3681) );
  OR3XL U5723 ( .A(input_previous_0[5]), .B(input_previous_0[6]), .C(n3635), 
        .Y(n3633) );
  OR3XL U5724 ( .A(input_previous_2[5]), .B(input_previous_2[6]), .C(n3731), 
        .Y(n3729) );
  OR3XL U5725 ( .A(output_previous_2[5]), .B(output_previous_2[6]), .C(n3827), 
        .Y(n3825) );
  OR3XL U5726 ( .A(input_previous_1[1]), .B(input_previous_1[2]), 
        .C(input_p1_times_b1_mul_componentxinput_A_inverted[0]), .Y(n3685) );
  OR3XL U5727 ( .A(input_previous_0[1]), .B(input_previous_0[2]), 
        .C(input_times_b0_mul_componentxinput_A_inverted[0]), .Y(n3637) );
  OR3XL U5728 ( .A(input_previous_2[1]), .B(input_previous_2[2]), 
        .C(input_p2_times_b2_mul_componentxinput_A_inverted[0]), .Y(n3733) );
  OR3XL U5729 ( .A(output_previous_2[1]), .B(output_previous_2[2]), 
        .C(output_p2_times_a2_mul_componentxinput_A_inverted[0]), .Y(n3829) );
  OR3XL U5730 ( .A(input_previous_1[3]), .B(input_previous_1[4]), .C(n3685), 
        .Y(n3683) );
  OR3XL U5731 ( .A(input_previous_0[3]), .B(input_previous_0[4]), .C(n3637), 
        .Y(n3635) );
  OR3XL U5732 ( .A(input_previous_2[3]), .B(input_previous_2[4]), .C(n3733), 
        .Y(n3731) );
  OR3XL U5733 ( .A(output_previous_2[3]), .B(output_previous_2[4]), .C(n3829), 
        .Y(n3827) );
  INVX1 U5734 ( .A(n4205), .Y(n373) );
  AOI22X1 U5735 ( .A0(n4203), 
        .A1(input_p1_times_b1_div_componentxoutput_sign_gated_prev), 
        .B0(n4204), .B1(n374), .Y(n4205) );
  XNOR2X1 U5736 ( .A(n124), .B(n333), .Y(n4204) );
  INVX1 U5737 ( .A(n4261), .Y(n375) );
  AOI22X1 U5738 ( .A0(n4259), 
        .A1(input_p2_times_b2_div_componentxoutput_sign_gated_prev), 
        .B0(n4260), .B1(n376), .Y(n4261) );
  XNOR2X1 U5739 ( .A(n128), .B(n324), .Y(n4260) );
  INVX1 U5740 ( .A(n4371), .Y(n377) );
  AOI22X1 U5741 ( .A0(n4369), 
        .A1(output_p2_times_a2_div_componentxoutput_sign_gated_prev), 
        .B0(n4370), .B1(n378), .Y(n4371) );
  XNOR2X1 U5742 ( .A(n116), .B(n351), .Y(n4370) );
  INVX1 U5743 ( .A(input_times_b0_div_componentxn27), .Y(n379) );
  AOI22X1 U5744 ( .A0(input_times_b0_div_componentxn24), 
        .A1(input_times_b0_div_componentxoutput_sign_gated_prev), 
        .B0(input_times_b0_div_componentxn25), .B1(n380), 
        .Y(input_times_b0_div_componentxn27) );
  XNOR2X1 U5745 ( .A(n120), .B(n342), .Y(input_times_b0_div_componentxn25) );
  BUFX3 U5746 ( .A(n4424), .Y(n180) );
  AOI22X1 U5747 ( .A0(input_previous_1[9]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[9]), 
        .B1(input_previous_1[17]), .Y(n4424) );
  XNOR2X1 U5748 ( .A(n3679), .B(input_previous_1[9]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[9]) );
  BUFX3 U5749 ( .A(n4477), .Y(n201) );
  AOI22X1 U5750 ( .A0(input_previous_2[9]), .A1(n142), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[9]), 
        .B1(input_previous_2[17]), .Y(n4477) );
  XNOR2X1 U5751 ( .A(n3727), .B(input_previous_2[9]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[9]) );
  BUFX3 U5752 ( .A(n4583), .Y(n243) );
  AOI22X1 U5753 ( .A0(output_previous_2[9]), .A1(n140), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[9]), 
        .B1(output_previous_2[17]), .Y(n4583) );
  XNOR2X1 U5754 ( .A(n3823), .B(output_previous_2[9]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[9]) );
  BUFX3 U5755 ( .A(input_times_b0_mul_componentxn73), .Y(n271) );
  AOI22X1 U5756 ( .A0(input_previous_0[9]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[9]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn73) );
  XNOR2X1 U5757 ( .A(n3631), .B(input_previous_0[9]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[9]) );
  OAI2BB1X1 U5758 ( 
        .A0N(input_p1_times_b1_div_componentxUDxshifted_substraction_result_0), 
        .A1N(n370), .B0(n1869), .Y(n1889) );
  AOI22X1 U5759 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_16), 
        .A1(n1870), .B0(input_p1_times_b1_div_componentxunsigned_A_17), 
        .B1(n1871), .Y(n1869) );
  NOR2BX1 U5760 ( .AN(input_p1_times_b1_div_componentxinput_A_inverted[17]), 
        .B(n190), .Y(input_p1_times_b1_div_componentxunsigned_A_17) );
  XOR2X1 U5761 ( .A(n3919), .B(n123), 
        .Y(input_p1_times_b1_div_componentxinput_A_inverted[17]) );
  OAI2BB1X1 U5762 ( 
        .A0N(input_p2_times_b2_div_componentxUDxshifted_substraction_result_0), 
        .A1N(n369), .B0(n1979), .Y(n1998) );
  AOI22X1 U5763 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_16), 
        .A1(n1980), .B0(input_p2_times_b2_div_componentxunsigned_A_17), 
        .B1(n1), .Y(n1979) );
  NOR2BX1 U5764 ( .AN(input_p2_times_b2_div_componentxinput_A_inverted[17]), 
        .B(n211), .Y(input_p2_times_b2_div_componentxunsigned_A_17) );
  XOR2X1 U5765 ( .A(n3962), .B(n127), 
        .Y(input_p2_times_b2_div_componentxinput_A_inverted[17]) );
  OAI2BB1X1 U5766 ( 
        .A0N(output_p2_times_a2_div_componentxUDxshifted_substraction_result_0), 
        .A1N(n368), .B0(n2198), .Y(n2217) );
  AOI22X1 U5767 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_16), 
        .A1(n2199), .B0(output_p2_times_a2_div_componentxunsigned_A_17), 
        .B1(n2090), .Y(n2198) );
  NOR2BX1 U5768 ( .AN(output_p2_times_a2_div_componentxinput_A_inverted[17]), 
        .B(n253), .Y(output_p2_times_a2_div_componentxunsigned_A_17) );
  XOR2X1 U5769 ( .A(n4048), .B(n115), 
        .Y(output_p2_times_a2_div_componentxinput_A_inverted[17]) );
  OAI2BB1X1 U5770 ( 
        .A0N(input_times_b0_div_componentxUDxshifted_substraction_result_0), 
        .A1N(n368), .B0(input_times_b0_div_componentxUDxinput_containerxn2), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn22) );
  AOI22X1 U5771 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_16), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), 
        .B0(input_times_b0_div_componentxunsigned_A_17), .B1(n1871), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn2) );
  NOR2BX1 U5772 ( .AN(input_times_b0_div_componentxinput_A_inverted[17]), 
        .B(n281), .Y(input_times_b0_div_componentxunsigned_A_17) );
  XOR2X1 U5773 ( .A(n3876), .B(n119), 
        .Y(input_times_b0_div_componentxinput_A_inverted[17]) );
  OAI2BB1X1 U5774 ( .A0N(n372), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_1), 
        .B0(n1887), .Y(n1905) );
  AOI22X1 U5775 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_0), 
        .A1(n1870), .B0(n857), .B1(n1871), .Y(n1887) );
  INVX1 U5776 ( .A(n4207), .Y(n857) );
  AOI22X1 U5777 ( .A0(n994), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[1]), .B1(n124), 
        .Y(n4207) );
  OAI2BB1X1 U5778 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_2), 
        .B0(n1886), .Y(n1904) );
  AOI22X1 U5779 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_1), 
        .A1(n1870), .B0(n858), .B1(n1871), .Y(n1886) );
  INVX1 U5780 ( .A(n4208), .Y(n858) );
  AOI22X1 U5781 ( .A0(n993), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[2]), .B1(n124), 
        .Y(n4208) );
  OAI2BB1X1 U5782 ( .A0N(n367), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_3), 
        .B0(n1885), .Y(n1903) );
  AOI22X1 U5783 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_2), 
        .A1(n1870), .B0(n859), .B1(n1871), .Y(n1885) );
  INVX1 U5784 ( .A(n4209), .Y(n859) );
  AOI22X1 U5785 ( .A0(n986), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[3]), .B1(n124), 
        .Y(n4209) );
  OAI2BB1X1 U5786 ( .A0N(n371), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_4), 
        .B0(n1884), .Y(n1902) );
  AOI22X1 U5787 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_3), 
        .A1(n1870), .B0(n860), .B1(n1871), .Y(n1884) );
  INVX1 U5788 ( .A(n4210), .Y(n860) );
  AOI22X1 U5789 ( .A0(n980), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[4]), .B1(n124), 
        .Y(n4210) );
  OAI2BB1X1 U5790 ( .A0N(n368), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_5), 
        .B0(n1883), .Y(n1901) );
  AOI22X1 U5791 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_4), 
        .A1(n1870), .B0(n861), .B1(n1871), .Y(n1883) );
  INVX1 U5792 ( .A(n4211), .Y(n861) );
  AOI22X1 U5793 ( .A0(n972), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[5]), .B1(n124), 
        .Y(n4211) );
  OAI2BB1X1 U5794 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_6), 
        .B0(n1882), .Y(n1900) );
  AOI22X1 U5795 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_5), 
        .A1(n1870), .B0(n862), .B1(n1871), .Y(n1882) );
  INVX1 U5796 ( .A(n4212), .Y(n862) );
  AOI22X1 U5797 ( .A0(n965), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[6]), .B1(n124), 
        .Y(n4212) );
  OAI2BB1X1 U5798 ( .A0N(n372), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_7), 
        .B0(n1881), .Y(n1899) );
  AOI22X1 U5799 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_6), 
        .A1(n1870), .B0(n863), .B1(n1871), .Y(n1881) );
  INVX1 U5800 ( .A(n4213), .Y(n863) );
  AOI22X1 U5801 ( .A0(n957), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[7]), .B1(n124), 
        .Y(n4213) );
  OAI2BB1X1 U5802 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_8), 
        .B0(n1880), .Y(n1898) );
  AOI22X1 U5803 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_7), 
        .A1(n1870), .B0(n864), .B1(n1871), .Y(n1880) );
  INVX1 U5804 ( .A(n4214), .Y(n864) );
  AOI22X1 U5805 ( .A0(n950), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[8]), .B1(n124), 
        .Y(n4214) );
  OAI2BB1X1 U5806 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_9), 
        .B0(n1879), .Y(n1897) );
  AOI22X1 U5807 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_8), 
        .A1(n1870), .B0(n865), .B1(n1871), .Y(n1879) );
  INVX1 U5808 ( .A(n4215), .Y(n865) );
  AOI22X1 U5809 ( .A0(n940), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[9]), .B1(n123), 
        .Y(n4215) );
  OAI2BB1X1 U5810 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_10), 
        .B0(n1878), .Y(n1896) );
  AOI22X1 U5811 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_9), 
        .A1(n1870), .B0(n866), .B1(n1871), .Y(n1878) );
  INVX1 U5812 ( .A(n4216), .Y(n866) );
  AOI22X1 U5813 ( .A0(n930), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[10]), .B1(n123), 
        .Y(n4216) );
  OAI2BB1X1 U5814 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_11), 
        .B0(n1877), .Y(n1895) );
  AOI22X1 U5815 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_10), 
        .A1(n1870), .B0(n867), .B1(n1871), .Y(n1877) );
  INVX1 U5816 ( .A(n4217), .Y(n867) );
  AOI22X1 U5817 ( .A0(n917), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[11]), .B1(n123), 
        .Y(n4217) );
  OAI2BB1X1 U5818 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_12), 
        .B0(n1876), .Y(n1894) );
  AOI22X1 U5819 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_11), 
        .A1(n1870), .B0(n868), .B1(n1871), .Y(n1876) );
  INVX1 U5820 ( .A(n4218), .Y(n868) );
  AOI22X1 U5821 ( .A0(n908), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[12]), .B1(n123), 
        .Y(n4218) );
  OAI2BB1X1 U5822 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_13), 
        .B0(n1875), .Y(n1893) );
  AOI22XL U5823 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_12), 
        .A1(n1870), .B0(n869), .B1(n1871), .Y(n1875) );
  INVX1 U5824 ( .A(n4219), .Y(n869) );
  AOI22X1 U5825 ( .A0(n899), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[13]), .B1(n123), 
        .Y(n4219) );
  OAI2BB1X1 U5826 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_14), 
        .B0(n1874), .Y(n1892) );
  AOI22XL U5827 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_13), 
        .A1(n1870), .B0(n870), .B1(n1871), .Y(n1874) );
  INVX1 U5828 ( .A(n4220), .Y(n870) );
  AOI22X1 U5829 ( .A0(n893), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[14]), .B1(n123), 
        .Y(n4220) );
  OAI2BB1X1 U5830 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_15), 
        .B0(n1873), .Y(n1891) );
  AOI22XL U5831 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_14), 
        .A1(n1870), .B0(n871), .B1(n1871), .Y(n1873) );
  INVX1 U5832 ( .A(n4221), .Y(n871) );
  AOI22X1 U5833 ( .A0(n884), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[15]), .B1(n123), 
        .Y(n4221) );
  OAI2BB1X1 U5834 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_16), 
        .B0(n1872), .Y(n1890) );
  AOI22XL U5835 ( 
        .A0(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_15), 
        .A1(n1870), .B0(n872), .B1(n1871), .Y(n1872) );
  INVX1 U5836 ( .A(n4222), .Y(n872) );
  AOI22X1 U5837 ( .A0(n876), .A1(n190), 
        .B0(input_p1_times_b1_div_componentxinput_A_inverted[16]), .B1(n123), 
        .Y(n4222) );
  OAI2BB1X1 U5838 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_1), 
        .B0(n1996), .Y(n2014) );
  AOI22X1 U5839 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_0), 
        .A1(n1980), .B0(n1016), .B1(n1), .Y(n1996) );
  INVX1 U5840 ( .A(n4263), .Y(n1016) );
  AOI22X1 U5841 ( .A0(n1153), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[1]), .B1(n128), 
        .Y(n4263) );
  OAI2BB1X1 U5842 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_2), 
        .B0(n1995), .Y(n2013) );
  AOI22X1 U5843 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_1), 
        .A1(n1980), .B0(n1017), .B1(n1), .Y(n1995) );
  INVX1 U5844 ( .A(n4264), .Y(n1017) );
  AOI22X1 U5845 ( .A0(n1152), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[2]), .B1(n128), 
        .Y(n4264) );
  OAI2BB1X1 U5846 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_3), 
        .B0(n1994), .Y(n2012) );
  AOI22X1 U5847 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_2), 
        .A1(n1980), .B0(n1018), .B1(n1), .Y(n1994) );
  INVX1 U5848 ( .A(n4265), .Y(n1018) );
  AOI22X1 U5849 ( .A0(n1145), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[3]), .B1(n128), 
        .Y(n4265) );
  OAI2BB1X1 U5850 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_4), 
        .B0(n1993), .Y(n2011) );
  AOI22X1 U5851 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_3), 
        .A1(n1980), .B0(n1019), .B1(n1), .Y(n1993) );
  INVX1 U5852 ( .A(n4266), .Y(n1019) );
  AOI22X1 U5853 ( .A0(n1139), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[4]), .B1(n128), 
        .Y(n4266) );
  OAI2BB1X1 U5854 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_5), 
        .B0(n1992), .Y(n2010) );
  AOI22X1 U5855 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_4), 
        .A1(n1980), .B0(n1020), .B1(n1), .Y(n1992) );
  INVX1 U5856 ( .A(n4267), .Y(n1020) );
  AOI22X1 U5857 ( .A0(n1131), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[5]), .B1(n128), 
        .Y(n4267) );
  OAI2BB1X1 U5858 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_6), 
        .B0(n1991), .Y(n2009) );
  AOI22X1 U5859 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_5), 
        .A1(n1980), .B0(n1021), .B1(n1), .Y(n1991) );
  INVX1 U5860 ( .A(n4268), .Y(n1021) );
  AOI22X1 U5861 ( .A0(n1124), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[6]), .B1(n128), 
        .Y(n4268) );
  OAI2BB1X1 U5862 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_7), 
        .B0(n1990), .Y(n2008) );
  AOI22X1 U5863 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_6), 
        .A1(n1980), .B0(n1022), .B1(n1), .Y(n1990) );
  INVX1 U5864 ( .A(n4269), .Y(n1022) );
  AOI22X1 U5865 ( .A0(n1116), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[7]), .B1(n128), 
        .Y(n4269) );
  OAI2BB1X1 U5866 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_8), 
        .B0(n1989), .Y(n2007) );
  AOI22X1 U5867 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_7), 
        .A1(n1980), .B0(n1023), .B1(n1), .Y(n1989) );
  INVX1 U5868 ( .A(n4270), .Y(n1023) );
  AOI22X1 U5869 ( .A0(n1109), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[8]), .B1(n128), 
        .Y(n4270) );
  OAI2BB1X1 U5870 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_9), 
        .B0(n1988), .Y(n2006) );
  AOI22X1 U5871 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_8), 
        .A1(n1980), .B0(n1024), .B1(n1), .Y(n1988) );
  INVX1 U5872 ( .A(n4271), .Y(n1024) );
  AOI22X1 U5873 ( .A0(n1099), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[9]), .B1(n127), 
        .Y(n4271) );
  OAI2BB1X1 U5874 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_10), 
        .B0(n1987), .Y(n2005) );
  AOI22X1 U5875 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_9), 
        .A1(n1980), .B0(n1025), .B1(n1), .Y(n1987) );
  INVX1 U5876 ( .A(n4272), .Y(n1025) );
  AOI22X1 U5877 ( .A0(n1089), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[10]), .B1(n127), 
        .Y(n4272) );
  OAI2BB1X1 U5878 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_11), 
        .B0(n1986), .Y(n2004) );
  AOI22X1 U5879 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_10), 
        .A1(n1980), .B0(n1026), .B1(n1), .Y(n1986) );
  INVX1 U5880 ( .A(n4273), .Y(n1026) );
  AOI22X1 U5881 ( .A0(n1076), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[11]), .B1(n127), 
        .Y(n4273) );
  OAI2BB1X1 U5882 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_12), 
        .B0(n1985), .Y(n2003) );
  AOI22X1 U5883 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_11), 
        .A1(n1980), .B0(n1027), .B1(n1), .Y(n1985) );
  INVX1 U5884 ( .A(n4274), .Y(n1027) );
  AOI22X1 U5885 ( .A0(n1067), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[12]), .B1(n127), 
        .Y(n4274) );
  OAI2BB1X1 U5886 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_13), 
        .B0(n1984), .Y(n2002) );
  AOI22XL U5887 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_12), 
        .A1(n1980), .B0(n1028), .B1(n1), .Y(n1984) );
  INVX1 U5888 ( .A(n4275), .Y(n1028) );
  AOI22X1 U5889 ( .A0(n1058), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[13]), .B1(n127), 
        .Y(n4275) );
  OAI2BB1X1 U5890 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_14), 
        .B0(n1983), .Y(n2001) );
  AOI22XL U5891 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_13), 
        .A1(n1980), .B0(n1029), .B1(n1), .Y(n1983) );
  INVX1 U5892 ( .A(n4276), .Y(n1029) );
  AOI22X1 U5893 ( .A0(n1052), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[14]), .B1(n127), 
        .Y(n4276) );
  OAI2BB1X1 U5894 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_15), 
        .B0(n1982), .Y(n2000) );
  AOI22XL U5895 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_14), 
        .A1(n1980), .B0(n1030), .B1(n1), .Y(n1982) );
  INVX1 U5896 ( .A(n4277), .Y(n1030) );
  AOI22X1 U5897 ( .A0(n1043), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[15]), .B1(n127), 
        .Y(n4277) );
  OAI2BB1X1 U5898 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_16), 
        .B0(n1981), .Y(n1999) );
  AOI22XL U5899 ( 
        .A0(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_15), 
        .A1(n1980), .B0(n1031), .B1(n1), .Y(n1981) );
  INVX1 U5900 ( .A(n4278), .Y(n1031) );
  AOI22X1 U5901 ( .A0(n1035), .A1(n211), 
        .B0(input_p2_times_b2_div_componentxinput_A_inverted[16]), .B1(n127), 
        .Y(n4278) );
  OAI2BB1X1 U5902 ( .A0N(n370), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_1), 
        .B0(n2215), .Y(n2233) );
  AOI22X1 U5903 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_0), 
        .A1(n2199), .B0(n539), .B1(n1871), .Y(n2215) );
  INVX1 U5904 ( .A(n4373), .Y(n539) );
  AOI22X1 U5905 ( .A0(n676), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[1]), .B1(n116), 
        .Y(n4373) );
  OAI2BB1X1 U5906 ( .A0N(n369), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_2), 
        .B0(n2214), .Y(n2232) );
  AOI22X1 U5907 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_1), 
        .A1(n2199), .B0(n540), .B1(n1), .Y(n2214) );
  INVX1 U5908 ( .A(n4374), .Y(n540) );
  AOI22X1 U5909 ( .A0(n675), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[2]), .B1(n116), 
        .Y(n4374) );
  OAI2BB1X1 U5910 ( .A0N(n367), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_3), 
        .B0(n2213), .Y(n2231) );
  AOI22X1 U5911 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_2), 
        .A1(n2199), .B0(n541), .B1(n2090), .Y(n2213) );
  INVX1 U5912 ( .A(n4375), .Y(n541) );
  AOI22X1 U5913 ( .A0(n668), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[3]), .B1(n116), 
        .Y(n4375) );
  OAI2BB1X1 U5914 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_4), 
        .B0(n2212), .Y(n2230) );
  AOI22X1 U5915 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_3), 
        .A1(n2199), .B0(n542), .B1(n1871), .Y(n2212) );
  INVX1 U5916 ( .A(n4376), .Y(n542) );
  AOI22X1 U5917 ( .A0(n662), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[4]), .B1(n116), 
        .Y(n4376) );
  OAI2BB1X1 U5918 ( .A0N(n370), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_5), 
        .B0(n2211), .Y(n2229) );
  AOI22X1 U5919 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_4), 
        .A1(n2199), .B0(n543), .B1(n1), .Y(n2211) );
  INVX1 U5920 ( .A(n4377), .Y(n543) );
  AOI22X1 U5921 ( .A0(n654), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[5]), .B1(n116), 
        .Y(n4377) );
  OAI2BB1X1 U5922 ( .A0N(n367), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_6), 
        .B0(n2210), .Y(n2228) );
  AOI22X1 U5923 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_5), 
        .A1(n2199), .B0(n544), .B1(n2090), .Y(n2210) );
  INVX1 U5924 ( .A(n4378), .Y(n544) );
  AOI22X1 U5925 ( .A0(n647), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[6]), .B1(n116), 
        .Y(n4378) );
  OAI2BB1X1 U5926 ( .A0N(n368), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_7), 
        .B0(n2209), .Y(n2227) );
  AOI22X1 U5927 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_6), 
        .A1(n2199), .B0(n545), .B1(n1871), .Y(n2209) );
  INVX1 U5928 ( .A(n4379), .Y(n545) );
  AOI22X1 U5929 ( .A0(n639), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[7]), .B1(n116), 
        .Y(n4379) );
  OAI2BB1X1 U5930 ( .A0N(n369), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_8), 
        .B0(n2208), .Y(n2226) );
  AOI22X1 U5931 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_7), 
        .A1(n2199), .B0(n546), .B1(n1), .Y(n2208) );
  INVX1 U5932 ( .A(n4380), .Y(n546) );
  AOI22X1 U5933 ( .A0(n632), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[8]), .B1(n116), 
        .Y(n4380) );
  OAI2BB1X1 U5934 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_9), 
        .B0(n2207), .Y(n2225) );
  AOI22X1 U5935 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_8), 
        .A1(n2199), .B0(n547), .B1(n2090), .Y(n2207) );
  INVX1 U5936 ( .A(n4381), .Y(n547) );
  AOI22X1 U5937 ( .A0(n622), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[9]), .B1(n115), 
        .Y(n4381) );
  OAI2BB1X1 U5938 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_10), 
        .B0(n2206), .Y(n2224) );
  AOI22X1 U5939 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_9), 
        .A1(n2199), .B0(n548), .B1(n1871), .Y(n2206) );
  INVX1 U5940 ( .A(n4382), .Y(n548) );
  AOI22X1 U5941 ( .A0(n612), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[10]), .B1(n115), 
        .Y(n4382) );
  OAI2BB1X1 U5942 ( .A0N(n370), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_11), 
        .B0(n2205), .Y(n2223) );
  AOI22X1 U5943 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_10), 
        .A1(n2199), .B0(n549), .B1(n1), .Y(n2205) );
  INVX1 U5944 ( .A(n4383), .Y(n549) );
  AOI22X1 U5945 ( .A0(n599), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[11]), .B1(n115), 
        .Y(n4383) );
  OAI2BB1X1 U5946 ( .A0N(n367), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_12), 
        .B0(n2204), .Y(n2222) );
  AOI22X1 U5947 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_11), 
        .A1(n2199), .B0(n550), .B1(n2090), .Y(n2204) );
  INVX1 U5948 ( .A(n4384), .Y(n550) );
  AOI22X1 U5949 ( .A0(n590), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[12]), .B1(n115), 
        .Y(n4384) );
  OAI2BB1X1 U5950 ( .A0N(n368), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_13), 
        .B0(n2203), .Y(n2221) );
  AOI22XL U5951 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_12), 
        .A1(n2199), .B0(n551), .B1(n1), .Y(n2203) );
  INVX1 U5952 ( .A(n4385), .Y(n551) );
  AOI22X1 U5953 ( .A0(n581), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[13]), .B1(n115), 
        .Y(n4385) );
  OAI2BB1X1 U5954 ( .A0N(n369), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_14), 
        .B0(n2202), .Y(n2220) );
  AOI22XL U5955 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_13), 
        .A1(n2199), .B0(n552), .B1(n2090), .Y(n2202) );
  INVX1 U5956 ( .A(n4386), .Y(n552) );
  AOI22X1 U5957 ( .A0(n575), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[14]), .B1(n115), 
        .Y(n4386) );
  OAI2BB1X1 U5958 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_15), 
        .B0(n2201), .Y(n2219) );
  AOI22XL U5959 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_14), 
        .A1(n2199), .B0(n553), .B1(n1871), .Y(n2201) );
  INVX1 U5960 ( .A(n4387), .Y(n553) );
  AOI22X1 U5961 ( .A0(n566), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[15]), .B1(n115), 
        .Y(n4387) );
  OAI2BB1X1 U5962 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_16), 
        .B0(n2200), .Y(n2218) );
  AOI22XL U5963 ( 
        .A0(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_15), 
        .A1(n2199), .B0(n554), .B1(n1), .Y(n2200) );
  INVX1 U5964 ( .A(n4388), .Y(n554) );
  AOI22X1 U5965 ( .A0(n558), .A1(n253), 
        .B0(output_p2_times_a2_div_componentxinput_A_inverted[16]), .B1(n115), 
        .Y(n4388) );
  OAI2BB1X1 U5966 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_1), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn20), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn38) );
  AOI22X1 U5967 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_0), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n698), 
        .B1(n1), .Y(input_times_b0_div_componentxUDxinput_containerxn20) );
  INVX1 U5968 ( .A(input_times_b0_div_componentxn29), .Y(n698) );
  AOI22X1 U5969 ( .A0(n835), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[1]), .B1(n120), 
        .Y(input_times_b0_div_componentxn29) );
  OAI2BB1X1 U5970 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_2), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn19), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn37) );
  AOI22X1 U5971 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_1), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n699), 
        .B1(n2090), .Y(input_times_b0_div_componentxUDxinput_containerxn19) );
  INVX1 U5972 ( .A(input_times_b0_div_componentxn30), .Y(n699) );
  AOI22X1 U5973 ( .A0(n834), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[2]), .B1(n120), 
        .Y(input_times_b0_div_componentxn30) );
  OAI2BB1X1 U5974 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_3), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn18), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn36) );
  AOI22X1 U5975 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_2), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n700), 
        .B1(n2090), .Y(input_times_b0_div_componentxUDxinput_containerxn18) );
  INVX1 U5976 ( .A(input_times_b0_div_componentxn31), .Y(n700) );
  AOI22X1 U5977 ( .A0(n827), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[3]), .B1(n120), 
        .Y(input_times_b0_div_componentxn31) );
  OAI2BB1X1 U5978 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_4), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn17), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn35) );
  AOI22X1 U5979 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_3), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n701), 
        .B1(n1871), .Y(input_times_b0_div_componentxUDxinput_containerxn17) );
  INVX1 U5980 ( .A(input_times_b0_div_componentxn32), .Y(n701) );
  AOI22X1 U5981 ( .A0(n821), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[4]), .B1(n120), 
        .Y(input_times_b0_div_componentxn32) );
  OAI2BB1X1 U5982 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_5), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn16), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn34) );
  AOI22X1 U5983 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_4), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n702), 
        .B1(n1), .Y(input_times_b0_div_componentxUDxinput_containerxn16) );
  INVX1 U5984 ( .A(input_times_b0_div_componentxn33), .Y(n702) );
  AOI22X1 U5985 ( .A0(n813), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[5]), .B1(n120), 
        .Y(input_times_b0_div_componentxn33) );
  OAI2BB1X1 U5986 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_6), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn15), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn33) );
  AOI22X1 U5987 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_5), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n703), 
        .B1(n2090), .Y(input_times_b0_div_componentxUDxinput_containerxn15) );
  INVX1 U5988 ( .A(input_times_b0_div_componentxn34), .Y(n703) );
  AOI22X1 U5989 ( .A0(n806), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[6]), .B1(n120), 
        .Y(input_times_b0_div_componentxn34) );
  OAI2BB1X1 U5990 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_7), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn14), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn32) );
  AOI22X1 U5991 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_6), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n704), 
        .B1(n1871), .Y(input_times_b0_div_componentxUDxinput_containerxn14) );
  INVX1 U5992 ( .A(input_times_b0_div_componentxn35), .Y(n704) );
  AOI22X1 U5993 ( .A0(n798), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[7]), .B1(n120), 
        .Y(input_times_b0_div_componentxn35) );
  OAI2BB1X1 U5994 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_8), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn13), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn31) );
  AOI22X1 U5995 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_7), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n705), 
        .B1(n1871), .Y(input_times_b0_div_componentxUDxinput_containerxn13) );
  INVX1 U5996 ( .A(input_times_b0_div_componentxn36), .Y(n705) );
  AOI22X1 U5997 ( .A0(n791), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[8]), .B1(n120), 
        .Y(input_times_b0_div_componentxn36) );
  OAI2BB1X1 U5998 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_9), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn12), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn30) );
  AOI22X1 U5999 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_8), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n706), 
        .B1(n1), .Y(input_times_b0_div_componentxUDxinput_containerxn12) );
  INVX1 U6000 ( .A(input_times_b0_div_componentxn37), .Y(n706) );
  AOI22X1 U6001 ( .A0(n781), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[9]), .B1(n119), 
        .Y(input_times_b0_div_componentxn37) );
  OAI2BB1X1 U6002 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_10), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn11), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn29) );
  AOI22X1 U6003 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_9), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n707), 
        .B1(n2090), .Y(input_times_b0_div_componentxUDxinput_containerxn11) );
  INVX1 U6004 ( .A(input_times_b0_div_componentxn38), .Y(n707) );
  AOI22X1 U6005 ( .A0(n771), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[10]), .B1(n119), 
        .Y(input_times_b0_div_componentxn38) );
  OAI2BB1X1 U6006 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_11), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn10), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn28) );
  AOI22X1 U6007 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_10), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n708), 
        .B1(n1), .Y(input_times_b0_div_componentxUDxinput_containerxn10) );
  INVX1 U6008 ( .A(input_times_b0_div_componentxn39), .Y(n708) );
  AOI22X1 U6009 ( .A0(n758), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[11]), .B1(n119), 
        .Y(input_times_b0_div_componentxn39) );
  OAI2BB1X1 U6010 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_12), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn9), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn27) );
  AOI22X1 U6011 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_11), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n709), 
        .B1(n1871), .Y(input_times_b0_div_componentxUDxinput_containerxn9) );
  INVX1 U6012 ( .A(input_times_b0_div_componentxn40), .Y(n709) );
  AOI22X1 U6013 ( .A0(n749), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[12]), .B1(n119), 
        .Y(input_times_b0_div_componentxn40) );
  OAI2BB1X1 U6014 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_13), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn8), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn26) );
  AOI22XL U6015 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_12), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n710), 
        .B1(n1871), .Y(input_times_b0_div_componentxUDxinput_containerxn8) );
  INVX1 U6016 ( .A(input_times_b0_div_componentxn41), .Y(n710) );
  AOI22X1 U6017 ( .A0(n740), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[13]), .B1(n119), 
        .Y(input_times_b0_div_componentxn41) );
  OAI2BB1X1 U6018 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_14), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn7), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn25) );
  AOI22XL U6019 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_13), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n711), 
        .B1(n1), .Y(input_times_b0_div_componentxUDxinput_containerxn7) );
  INVX1 U6020 ( .A(input_times_b0_div_componentxn42), .Y(n711) );
  AOI22X1 U6021 ( .A0(n734), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[14]), .B1(n119), 
        .Y(input_times_b0_div_componentxn42) );
  OAI2BB1X1 U6022 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_15), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn6), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn24) );
  AOI22XL U6023 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_14), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n712), 
        .B1(n2090), .Y(input_times_b0_div_componentxUDxinput_containerxn6) );
  INVX1 U6024 ( .A(input_times_b0_div_componentxn43), .Y(n712) );
  AOI22X1 U6025 ( .A0(n725), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[15]), .B1(n119), 
        .Y(input_times_b0_div_componentxn43) );
  OAI2BB1X1 U6026 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_16), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn5), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn23) );
  AOI22XL U6027 ( 
        .A0(input_times_b0_div_componentxUDxinput_containerxparallel_out_15), 
        .A1(input_times_b0_div_componentxUDxinput_containerxn3), .B0(n713), 
        .B1(n2090), .Y(input_times_b0_div_componentxUDxinput_containerxn5) );
  INVX1 U6028 ( .A(input_times_b0_div_componentxn44), .Y(n713) );
  AOI22X1 U6029 ( .A0(n717), .A1(n281), 
        .B0(input_times_b0_div_componentxinput_A_inverted[16]), .B1(n119), 
        .Y(input_times_b0_div_componentxn44) );
  OAI2BB1X1 U6030 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_0), 
        .B0(n1888), .Y(n1906) );
  NAND2XL U6031 ( .A(n856), .B(n1871), .Y(n1888) );
  INVX1 U6032 ( .A(n4206), .Y(n856) );
  AOI22X1 U6033 ( .A0(n995), .A1(n190), .B0(n995), .B1(n124), .Y(n4206) );
  OAI2BB1X1 U6034 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_0), 
        .B0(n1997), .Y(n2015) );
  NAND2XL U6035 ( .A(n1015), .B(n1), .Y(n1997) );
  INVX1 U6036 ( .A(n4262), .Y(n1015) );
  AOI22X1 U6037 ( .A0(n1154), .A1(n211), .B0(n1154), .B1(n128), .Y(n4262) );
  OAI2BB1X1 U6038 ( .A0N(n367), 
        .A1N(output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_0), 
        .B0(n2216), .Y(n2234) );
  NAND2XL U6039 ( .A(n538), .B(n1871), .Y(n2216) );
  INVX1 U6040 ( .A(n4372), .Y(n538) );
  AOI22X1 U6041 ( .A0(n677), .A1(n253), .B0(n677), .B1(n116), .Y(n4372) );
  OAI2BB1X1 U6042 ( .A0N(n368), 
        .A1N(input_times_b0_div_componentxUDxinput_containerxparallel_out_0), 
        .B0(input_times_b0_div_componentxUDxinput_containerxn21), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn40) );
  NAND2XL U6043 ( .A(n697), .B(n1), 
        .Y(input_times_b0_div_componentxUDxinput_containerxn21) );
  INVX1 U6044 ( .A(input_times_b0_div_componentxn28), .Y(n697) );
  AOI22X1 U6045 ( .A0(n836), .A1(n281), .B0(n836), .B1(n120), 
        .Y(input_times_b0_div_componentxn28) );
  AOI22X1 U6046 ( .A0(input_previous_2[11]), .A1(n141), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[11]), 
        .B1(input_previous_2[17]), .Y(n4491) );
  XOR2X1 U6047 ( .A(n3740), .B(input_previous_2[11]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[11]) );
  AOI22X1 U6048 ( .A0(output_previous_2[11]), .A1(n139), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[11]), 
        .B1(output_previous_2[17]), .Y(n4597) );
  XOR2X1 U6049 ( .A(n3836), .B(output_previous_2[11]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[11]) );
  AOI22X1 U6050 ( .A0(input_previous_2[12]), .A1(n141), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[12]), 
        .B1(input_previous_2[17]), .Y(n4490) );
  XOR2X1 U6051 ( .A(n3741), .B(input_previous_2[12]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[12]) );
  OR2X2 U6052 ( .A(n3740), .B(input_previous_2[11]), .Y(n3741) );
  AOI22X1 U6053 ( .A0(output_previous_2[12]), .A1(n139), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[12]), 
        .B1(output_previous_2[17]), .Y(n4596) );
  XOR2X1 U6054 ( .A(n3837), .B(output_previous_2[12]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[12]) );
  OR2X2 U6055 ( .A(n3836), .B(output_previous_2[11]), .Y(n3837) );
  AOI22X1 U6056 ( .A0(input_previous_1[13]), .A1(n143), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[13]), 
        .B1(input_previous_1[17]), .Y(n4436) );
  XOR2X1 U6057 ( .A(n3690), .B(input_previous_1[13]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[13]) );
  AOI22X1 U6058 ( .A0(input_previous_2[13]), .A1(n141), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[13]), 
        .B1(input_previous_2[17]), .Y(n4489) );
  XOR2X1 U6059 ( .A(n3738), .B(input_previous_2[13]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[13]) );
  AOI22X1 U6060 ( .A0(output_previous_2[13]), .A1(n139), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[13]), 
        .B1(output_previous_2[17]), .Y(n4595) );
  XOR2X1 U6061 ( .A(n3834), .B(output_previous_2[13]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[13]) );
  AOI22X1 U6062 ( .A0(input_previous_0[13]), .A1(n131), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[13]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn85) );
  XOR2X1 U6063 ( .A(n3642), .B(input_previous_0[13]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[13]) );
  AOI22X1 U6064 ( .A0(input_previous_1[14]), .A1(n143), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[14]), 
        .B1(input_previous_1[17]), .Y(n4435) );
  XOR2X1 U6065 ( .A(n3691), .B(input_previous_1[14]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[14]) );
  OR2X2 U6066 ( .A(input_previous_1[13]), .B(n3690), .Y(n3691) );
  AOI22X1 U6067 ( .A0(input_previous_2[14]), .A1(n141), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[14]), 
        .B1(input_previous_2[17]), .Y(n4488) );
  XOR2X1 U6068 ( .A(n3739), .B(input_previous_2[14]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[14]) );
  OR2X2 U6069 ( .A(input_previous_2[13]), .B(n3738), .Y(n3739) );
  AOI22X1 U6070 ( .A0(output_previous_2[14]), .A1(n139), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[14]), 
        .B1(output_previous_2[17]), .Y(n4594) );
  XOR2X1 U6071 ( .A(n3835), .B(output_previous_2[14]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[14]) );
  OR2X2 U6072 ( .A(output_previous_2[13]), .B(n3834), .Y(n3835) );
  AOI22X1 U6073 ( .A0(input_previous_0[14]), .A1(n131), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[14]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn84) );
  XOR2X1 U6074 ( .A(n3643), .B(input_previous_0[14]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[14]) );
  OR2X2 U6075 ( .A(input_previous_0[13]), .B(n3642), .Y(n3643) );
  AOI22X1 U6076 ( .A0(input_previous_2[15]), .A1(n141), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[15]), 
        .B1(input_previous_2[17]), .Y(n4487) );
  XNOR2X1 U6077 ( .A(n3737), .B(input_previous_2[15]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[15]) );
  AOI22X1 U6078 ( .A0(output_previous_2[15]), .A1(n139), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[15]), 
        .B1(output_previous_2[17]), .Y(n4593) );
  XNOR2X1 U6079 ( .A(n3833), .B(output_previous_2[15]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[15]) );
  NOR3X1 U6080 ( .A(input_previous_1[13]), .B(input_previous_1[14]), .C(n3690), 
        .Y(n3689) );
  NOR3X1 U6081 ( .A(input_previous_0[13]), .B(input_previous_0[14]), .C(n3642), 
        .Y(n3641) );
  NOR3X1 U6082 ( .A(input_previous_2[13]), .B(input_previous_2[14]), .C(n3738), 
        .Y(n3737) );
  NOR3X1 U6083 ( .A(output_previous_2[13]), .B(output_previous_2[14]), 
        .C(n3834), .Y(n3833) );
  BUFX3 U6084 ( .A(n4429), .Y(n185) );
  AOI22X1 U6085 ( .A0(input_previous_1[4]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[4]), 
        .B1(input_previous_1[17]), .Y(n4429) );
  XOR2X1 U6086 ( .A(n3684), .B(input_previous_1[4]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[4]) );
  OR2X2 U6087 ( .A(input_previous_1[3]), .B(n3685), .Y(n3684) );
  BUFX3 U6088 ( .A(input_times_b0_mul_componentxn78), .Y(n276) );
  AOI22X1 U6089 ( .A0(input_previous_0[4]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[4]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn78) );
  XOR2X1 U6090 ( .A(n3636), .B(input_previous_0[4]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[4]) );
  OR2X2 U6091 ( .A(input_previous_0[3]), .B(n3637), .Y(n3636) );
  NAND3BX1 U6092 ( .AN(input_previous_2[10]), .B(n1283), .C(n3727), .Y(n3740)
         );
  NAND3BX1 U6093 ( .AN(output_previous_2[10]), .B(n1282), .C(n3823), .Y(n3836)
         );
  OR3XL U6094 ( .A(input_previous_1[11]), .B(input_previous_1[12]), .C(n3692), 
        .Y(n3690) );
  OR3XL U6095 ( .A(input_previous_0[11]), .B(input_previous_0[12]), .C(n3644), 
        .Y(n3642) );
  OR3XL U6096 ( .A(input_previous_2[11]), .B(input_previous_2[12]), .C(n3740), 
        .Y(n3738) );
  OR3XL U6097 ( .A(output_previous_2[11]), .B(output_previous_2[12]), 
        .C(n3836), .Y(n3834) );
  BUFX3 U6098 ( .A(n4440), .Y(n189) );
  AOI22X1 U6099 ( .A0(input_p1_times_b1_mul_componentxinput_A_inverted[0]), 
        .A1(n143), .B0(input_p1_times_b1_mul_componentxinput_A_inverted[0]), 
        .B1(input_previous_1[17]), .Y(n4440) );
  BUFX3 U6100 ( .A(n4493), .Y(n210) );
  AOI22X1 U6101 ( .A0(input_p2_times_b2_mul_componentxinput_A_inverted[0]), 
        .A1(n141), .B0(input_p2_times_b2_mul_componentxinput_A_inverted[0]), 
        .B1(input_previous_2[17]), .Y(n4493) );
  BUFX3 U6102 ( .A(n4599), .Y(n252) );
  AOI22X1 U6103 ( .A0(output_p2_times_a2_mul_componentxinput_A_inverted[0]), 
        .A1(n139), .B0(output_p2_times_a2_mul_componentxinput_A_inverted[0]), 
        .B1(output_previous_2[17]), .Y(n4599) );
  BUFX3 U6104 ( .A(input_times_b0_mul_componentxn89), .Y(n280) );
  AOI22X1 U6105 ( .A0(input_times_b0_mul_componentxinput_A_inverted[0]), 
        .A1(n131), .B0(input_times_b0_mul_componentxinput_A_inverted[0]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn89) );
  BUFX3 U6106 ( .A(n4432), .Y(n188) );
  AOI22X1 U6107 ( .A0(input_previous_1[1]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[1]), 
        .B1(input_previous_1[17]), .Y(n4432) );
  XOR2X1 U6108 ( .A(input_previous_1[1]), 
        .B(input_p1_times_b1_mul_componentxinput_A_inverted[0]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[1]) );
  BUFX3 U6109 ( .A(n4485), .Y(n209) );
  AOI22X1 U6110 ( .A0(input_previous_2[1]), .A1(n141), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[1]), 
        .B1(input_previous_2[17]), .Y(n4485) );
  XOR2X1 U6111 ( .A(input_previous_2[1]), 
        .B(input_p2_times_b2_mul_componentxinput_A_inverted[0]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[1]) );
  BUFX3 U6112 ( .A(n4591), .Y(n251) );
  AOI22X1 U6113 ( .A0(output_previous_2[1]), .A1(n139), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[1]), 
        .B1(output_previous_2[17]), .Y(n4591) );
  XOR2X1 U6114 ( .A(output_previous_2[1]), 
        .B(output_p2_times_a2_mul_componentxinput_A_inverted[0]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[1]) );
  BUFX3 U6115 ( .A(input_times_b0_mul_componentxn81), .Y(n279) );
  AOI22X1 U6116 ( .A0(input_previous_0[1]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[1]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn81) );
  XOR2X1 U6117 ( .A(input_previous_0[1]), 
        .B(input_times_b0_mul_componentxinput_A_inverted[0]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[1]) );
  BUFX3 U6118 ( .A(n4431), .Y(n187) );
  AOI22X1 U6119 ( .A0(input_previous_1[2]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[2]), 
        .B1(input_previous_1[17]), .Y(n4431) );
  XNOR2X1 U6120 ( .A(input_previous_1[2]), .B(n3686), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[2]) );
  NOR2X1 U6121 ( .A(input_p1_times_b1_mul_componentxinput_A_inverted[0]), 
        .B(input_previous_1[1]), .Y(n3686) );
  BUFX3 U6122 ( .A(n4484), .Y(n208) );
  AOI22X1 U6123 ( .A0(input_previous_2[2]), .A1(n142), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[2]), 
        .B1(input_previous_2[17]), .Y(n4484) );
  XNOR2X1 U6124 ( .A(input_previous_2[2]), .B(n3734), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[2]) );
  NOR2X1 U6125 ( .A(input_p2_times_b2_mul_componentxinput_A_inverted[0]), 
        .B(input_previous_2[1]), .Y(n3734) );
  BUFX3 U6126 ( .A(n4590), .Y(n250) );
  AOI22X1 U6127 ( .A0(output_previous_2[2]), .A1(n140), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[2]), 
        .B1(output_previous_2[17]), .Y(n4590) );
  XNOR2X1 U6128 ( .A(output_previous_2[2]), .B(n3830), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[2]) );
  NOR2X1 U6129 ( .A(output_p2_times_a2_mul_componentxinput_A_inverted[0]), 
        .B(output_previous_2[1]), .Y(n3830) );
  BUFX3 U6130 ( .A(input_times_b0_mul_componentxn80), .Y(n278) );
  AOI22X1 U6131 ( .A0(input_previous_0[2]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[2]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn80) );
  XNOR2X1 U6132 ( .A(input_previous_0[2]), .B(n3638), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[2]) );
  NOR2X1 U6133 ( .A(input_times_b0_mul_componentxinput_A_inverted[0]), 
        .B(input_previous_0[1]), .Y(n3638) );
  BUFX3 U6134 ( .A(n4430), .Y(n186) );
  AOI22X1 U6135 ( .A0(input_previous_1[3]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[3]), 
        .B1(input_previous_1[17]), .Y(n4430) );
  XOR2X1 U6136 ( .A(n3685), .B(input_previous_1[3]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[3]) );
  BUFX3 U6137 ( .A(input_times_b0_mul_componentxn79), .Y(n277) );
  AOI22X1 U6138 ( .A0(input_previous_0[3]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[3]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn79) );
  XOR2X1 U6139 ( .A(n3637), .B(input_previous_0[3]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[3]) );
  BUFX3 U6140 ( .A(n4428), .Y(n184) );
  AOI22X1 U6141 ( .A0(input_previous_1[5]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[5]), 
        .B1(input_previous_1[17]), .Y(n4428) );
  XOR2X1 U6142 ( .A(n3683), .B(input_previous_1[5]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[5]) );
  BUFX3 U6143 ( .A(n4481), .Y(n205) );
  AOI22X1 U6144 ( .A0(input_previous_2[5]), .A1(n142), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[5]), 
        .B1(input_previous_2[17]), .Y(n4481) );
  XOR2X1 U6145 ( .A(n3731), .B(input_previous_2[5]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[5]) );
  BUFX3 U6146 ( .A(n4587), .Y(n247) );
  AOI22X1 U6147 ( .A0(output_previous_2[5]), .A1(n140), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[5]), 
        .B1(output_previous_2[17]), .Y(n4587) );
  XOR2X1 U6148 ( .A(n3827), .B(output_previous_2[5]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[5]) );
  BUFX3 U6149 ( .A(input_times_b0_mul_componentxn77), .Y(n275) );
  AOI22X1 U6150 ( .A0(input_previous_0[5]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[5]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn77) );
  XOR2X1 U6151 ( .A(n3635), .B(input_previous_0[5]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[5]) );
  BUFX3 U6152 ( .A(n4427), .Y(n183) );
  AOI22X1 U6153 ( .A0(input_previous_1[6]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[6]), 
        .B1(input_previous_1[17]), .Y(n4427) );
  XOR2X1 U6154 ( .A(n3682), .B(input_previous_1[6]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[6]) );
  OR2X2 U6155 ( .A(input_previous_1[5]), .B(n3683), .Y(n3682) );
  BUFX3 U6156 ( .A(n4480), .Y(n204) );
  AOI22X1 U6157 ( .A0(input_previous_2[6]), .A1(n142), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[6]), 
        .B1(input_previous_2[17]), .Y(n4480) );
  XOR2X1 U6158 ( .A(n3730), .B(input_previous_2[6]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[6]) );
  OR2X2 U6159 ( .A(input_previous_2[5]), .B(n3731), .Y(n3730) );
  BUFX3 U6160 ( .A(n4586), .Y(n246) );
  AOI22X1 U6161 ( .A0(output_previous_2[6]), .A1(n140), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[6]), 
        .B1(output_previous_2[17]), .Y(n4586) );
  XOR2X1 U6162 ( .A(n3826), .B(output_previous_2[6]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[6]) );
  OR2X2 U6163 ( .A(output_previous_2[5]), .B(n3827), .Y(n3826) );
  BUFX3 U6164 ( .A(input_times_b0_mul_componentxn76), .Y(n274) );
  AOI22X1 U6165 ( .A0(input_previous_0[6]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[6]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn76) );
  XOR2X1 U6166 ( .A(n3634), .B(input_previous_0[6]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[6]) );
  OR2X2 U6167 ( .A(input_previous_0[5]), .B(n3635), .Y(n3634) );
  BUFX3 U6168 ( .A(n4426), .Y(n182) );
  AOI22X1 U6169 ( .A0(input_previous_1[7]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[7]), 
        .B1(input_previous_1[17]), .Y(n4426) );
  XOR2X1 U6170 ( .A(n3681), .B(input_previous_1[7]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[7]) );
  BUFX3 U6171 ( .A(n4479), .Y(n203) );
  AOI22X1 U6172 ( .A0(input_previous_2[7]), .A1(n142), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[7]), 
        .B1(input_previous_2[17]), .Y(n4479) );
  XOR2X1 U6173 ( .A(n3729), .B(input_previous_2[7]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[7]) );
  BUFX3 U6174 ( .A(n4585), .Y(n245) );
  AOI22X1 U6175 ( .A0(output_previous_2[7]), .A1(n140), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[7]), 
        .B1(output_previous_2[17]), .Y(n4585) );
  XOR2X1 U6176 ( .A(n3825), .B(output_previous_2[7]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[7]) );
  BUFX3 U6177 ( .A(input_times_b0_mul_componentxn75), .Y(n273) );
  AOI22X1 U6178 ( .A0(input_previous_0[7]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[7]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn75) );
  XOR2X1 U6179 ( .A(n3633), .B(input_previous_0[7]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[7]) );
  AOI22X1 U6180 ( .A0(input_previous_1[15]), .A1(n143), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[15]), 
        .B1(input_previous_1[17]), .Y(n4434) );
  XNOR2X1 U6181 ( .A(n3689), .B(input_previous_1[15]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[15]) );
  AOI22X1 U6182 ( .A0(input_previous_0[15]), .A1(n131), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[15]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn83) );
  XNOR2X1 U6183 ( .A(n3641), .B(input_previous_0[15]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[15]) );
  INVX1 U6184 ( .A(input_previous_1[17]), .Y(n254) );
  INVX1 U6185 ( .A(input_previous_2[17]), .Y(n255) );
  INVX1 U6186 ( .A(output_previous_2[17]), .Y(n256) );
  INVX1 U6187 ( .A(input_previous_0[17]), .Y(n282) );
  BUFX3 U6188 ( .A(n4478), .Y(n202) );
  AOI22X1 U6189 ( .A0(input_previous_2[8]), .A1(n142), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[8]), 
        .B1(input_previous_2[17]), .Y(n4478) );
  XOR2X1 U6190 ( .A(n3728), .B(input_previous_2[8]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[8]) );
  OR2X2 U6191 ( .A(input_previous_2[7]), .B(n3729), .Y(n3728) );
  BUFX3 U6192 ( .A(n4584), .Y(n244) );
  AOI22X1 U6193 ( .A0(output_previous_2[8]), .A1(n140), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[8]), 
        .B1(output_previous_2[17]), .Y(n4584) );
  XOR2X1 U6194 ( .A(n3824), .B(output_previous_2[8]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[8]) );
  OR2X2 U6195 ( .A(output_previous_2[7]), .B(n3825), .Y(n3824) );
  BUFX3 U6196 ( .A(n4483), .Y(n207) );
  AOI22X1 U6197 ( .A0(input_previous_2[3]), .A1(n142), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[3]), 
        .B1(input_previous_2[17]), .Y(n4483) );
  XOR2X1 U6198 ( .A(n3733), .B(input_previous_2[3]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[3]) );
  BUFX3 U6199 ( .A(n4589), .Y(n249) );
  AOI22X1 U6200 ( .A0(output_previous_2[3]), .A1(n140), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[3]), 
        .B1(output_previous_2[17]), .Y(n4589) );
  XOR2X1 U6201 ( .A(n3829), .B(output_previous_2[3]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[3]) );
  AOI22X1 U6202 ( .A0(input_previous_1[12]), .A1(n143), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[12]), 
        .B1(input_previous_1[17]), .Y(n4437) );
  XOR2X1 U6203 ( .A(n3693), .B(input_previous_1[12]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[12]) );
  OR2X2 U6204 ( .A(n3692), .B(input_previous_1[11]), .Y(n3693) );
  AOI22X1 U6205 ( .A0(input_previous_0[12]), .A1(n131), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[12]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn86) );
  XOR2X1 U6206 ( .A(n3645), .B(input_previous_0[12]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[12]) );
  OR2X2 U6207 ( .A(n3644), .B(input_previous_0[11]), .Y(n3645) );
  BUFX3 U6208 ( .A(n4425), .Y(n181) );
  AOI22X1 U6209 ( .A0(input_previous_1[8]), .A1(n144), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[8]), 
        .B1(input_previous_1[17]), .Y(n4425) );
  XOR2X1 U6210 ( .A(n3680), .B(input_previous_1[8]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[8]) );
  OR2X2 U6211 ( .A(input_previous_1[7]), .B(n3681), .Y(n3680) );
  BUFX3 U6212 ( .A(input_times_b0_mul_componentxn74), .Y(n272) );
  AOI22X1 U6213 ( .A0(input_previous_0[8]), .A1(n132), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[8]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn74) );
  XOR2X1 U6214 ( .A(n3632), .B(input_previous_0[8]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[8]) );
  OR2X2 U6215 ( .A(input_previous_0[7]), .B(n3633), .Y(n3632) );
  BUFX3 U6216 ( .A(n4482), .Y(n206) );
  AOI22X1 U6217 ( .A0(input_previous_2[4]), .A1(n142), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[4]), 
        .B1(input_previous_2[17]), .Y(n4482) );
  XOR2X1 U6218 ( .A(n3732), .B(input_previous_2[4]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[4]) );
  OR2X2 U6219 ( .A(input_previous_2[3]), .B(n3733), .Y(n3732) );
  BUFX3 U6220 ( .A(n4588), .Y(n248) );
  AOI22X1 U6221 ( .A0(output_previous_2[4]), .A1(n140), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[4]), 
        .B1(output_previous_2[17]), .Y(n4588) );
  XOR2X1 U6222 ( .A(n3828), .B(output_previous_2[4]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[4]) );
  OR2X2 U6223 ( .A(output_previous_2[3]), .B(n3829), .Y(n3828) );
  AOI22X1 U6224 ( .A0(input_previous_1[16]), .A1(n143), 
        .B0(input_p1_times_b1_mul_componentxinput_A_inverted[16]), 
        .B1(input_previous_1[17]), .Y(n4433) );
  XNOR2X1 U6225 ( .A(n3688), .B(input_previous_1[16]), 
        .Y(input_p1_times_b1_mul_componentxinput_A_inverted[16]) );
  AOI22X1 U6226 ( .A0(input_previous_2[16]), .A1(n141), 
        .B0(input_p2_times_b2_mul_componentxinput_A_inverted[16]), 
        .B1(input_previous_2[17]), .Y(n4486) );
  XNOR2X1 U6227 ( .A(n3736), .B(input_previous_2[16]), 
        .Y(input_p2_times_b2_mul_componentxinput_A_inverted[16]) );
  AOI22X1 U6228 ( .A0(output_previous_2[16]), .A1(n139), 
        .B0(output_p2_times_a2_mul_componentxinput_A_inverted[16]), 
        .B1(output_previous_2[17]), .Y(n4592) );
  XNOR2X1 U6229 ( .A(n3832), .B(output_previous_2[16]), 
        .Y(output_p2_times_a2_mul_componentxinput_A_inverted[16]) );
  AOI22X1 U6230 ( .A0(input_previous_0[16]), .A1(n131), 
        .B0(input_times_b0_mul_componentxinput_A_inverted[16]), 
        .B1(input_previous_0[17]), .Y(input_times_b0_mul_componentxn82) );
  XNOR2X1 U6231 ( .A(n3640), .B(input_previous_0[16]), 
        .Y(input_times_b0_mul_componentxinput_A_inverted[16]) );
  NOR2BX1 U6232 ( .AN(n3689), .B(input_previous_1[15]), .Y(n3688) );
  NOR2BX1 U6233 ( .AN(n3641), .B(input_previous_0[15]), .Y(n3640) );
  NOR2BX1 U6234 ( .AN(n3737), .B(input_previous_2[15]), .Y(n3736) );
  NOR2BX1 U6235 ( .AN(n3833), .B(output_previous_2[15]), .Y(n3832) );
  INVX1 U6236 ( .A(input_previous_1[9]), .Y(n1293) );
  INVX1 U6237 ( .A(input_previous_0[9]), .Y(n1191) );
  NAND2BX1 U6238 ( .AN(input_previous_1[16]), .B(n3688), .Y(n3687) );
  NAND2BX1 U6239 ( .AN(input_previous_0[16]), .B(n3640), .Y(n3639) );
  NAND2BX1 U6240 ( .AN(input_previous_2[16]), .B(n3736), .Y(n3735) );
  NAND2BX1 U6241 ( .AN(output_previous_2[16]), .B(n3832), .Y(n3831) );
  INVX1 U6242 ( .A(input_previous_2[9]), .Y(n1283) );
  INVX1 U6243 ( .A(output_previous_2[9]), .Y(n1282) );
  OAI2BB2X1 U6244 ( .B0(n1214), .B1(n1260), .A0N(output_previous_2[7]), 
        .A1N(n320), .Y(n4662) );
  INVX1 U6245 ( .A(\output_signal[7] ), .Y(n1214) );
  OAI2BB2X1 U6246 ( .B0(n1218), .B1(n321), .A0N(output_previous_2[5]), 
        .A1N(n320), .Y(n4660) );
  INVX1 U6247 ( .A(\output_signal[5] ), .Y(n1218) );
  OAI2BB2X1 U6248 ( .B0(n1216), .B1(n1260), .A0N(output_previous_2[6]), 
        .A1N(n320), .Y(n4661) );
  INVX1 U6249 ( .A(\output_signal[6] ), .Y(n1216) );
  OAI2BB2X1 U6250 ( .B0(n1202), .B1(n1260), .A0N(output_previous_2[15]), 
        .A1N(n319), .Y(n4670) );
  INVX1 U6251 ( .A(output_previous_1[15]), .Y(n1202) );
  OAI2BB2X1 U6252 ( .B0(n1201), .B1(n320), .A0N(output_previous_2[14]), 
        .A1N(n319), .Y(n4669) );
  INVX1 U6253 ( .A(output_previous_1[14]), .Y(n1201) );
  OAI2BB2X1 U6254 ( .B0(n1200), .B1(n319), .A0N(output_previous_2[13]), 
        .A1N(n319), .Y(n4668) );
  INVX1 U6255 ( .A(output_previous_1[13]), .Y(n1200) );
  OAI2BB2X1 U6256 ( .B0(n1204), .B1(n1260), .A0N(output_previous_2[16]), 
        .A1N(n319), .Y(n4671) );
  INVX1 U6257 ( .A(output_previous_1[16]), .Y(n1204) );
  OAI2BB2X1 U6258 ( .B0(n1224), .B1(n1260), .A0N(output_previous_2[2]), 
        .A1N(n320), .Y(n4657) );
  INVX1 U6259 ( .A(\output_signal[2] ), .Y(n1224) );
  OAI2BB2X1 U6260 ( .B0(n1222), .B1(n319), .A0N(output_previous_2[3]), 
        .A1N(n320), .Y(n4658) );
  INVX1 U6261 ( .A(\output_signal[3] ), .Y(n1222) );
  OAI2BB2X1 U6262 ( .B0(n1220), .B1(n1260), .A0N(output_previous_2[4]), 
        .A1N(n320), .Y(n4659) );
  INVX1 U6263 ( .A(\output_signal[4] ), .Y(n1220) );
  OAI2BB2X1 U6264 ( .B0(n1206), .B1(n319), .A0N(output_previous_2[11]), 
        .A1N(n320), .Y(n4666) );
  INVX1 U6265 ( .A(output_previous_1[11]), .Y(n1206) );
  OAI2BB2X1 U6266 ( .B0(n1208), .B1(n1260), .A0N(output_previous_2[10]), 
        .A1N(n320), .Y(n4665) );
  INVX1 U6267 ( .A(output_previous_1[10]), .Y(n1208) );
  OAI2BB2X1 U6268 ( .B0(n1210), .B1(n321), .A0N(output_previous_2[9]), 
        .A1N(n320), .Y(n4664) );
  OAI2BB2X1 U6269 ( .B0(n1199), .B1(n1260), .A0N(output_previous_2[12]), 
        .A1N(n320), .Y(n4667) );
  INVX1 U6270 ( .A(output_previous_1[12]), .Y(n1199) );
  AOI32X1 U6271 ( .A0(n846), 
        .A1(input_times_b0_div_componentxUDxactually_substractsxn18), 
        .A2(input_times_b0_div_componentxUDxcentral_parallel_output_0), 
        .B0(input_times_b0_div_componentxUDxsub_ready_negative_divisor[1]), 
        .B1(input_times_b0_div_componentxUDxcentral_parallel_output_1), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn16) );
  AOI32X1 U6272 ( .A0(n1005), .A1(n1650), 
        .A2(input_p1_times_b1_div_componentxUDxcentral_parallel_output_0), 
        .B0(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[1]), 
        .B1(input_p1_times_b1_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1648) );
  AOI32X1 U6273 ( .A0(n1164), .A1(n1682), 
        .A2(input_p2_times_b2_div_componentxUDxcentral_parallel_output_0), 
        .B0(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[1]), 
        .B1(input_p2_times_b2_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1680) );
  AOI32X1 U6274 ( .A0(n528), .A1(n1714), 
        .A2(output_p1_times_a1_div_componentxUDxcentral_parallel_output_0), 
        .B0(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[1]), 
        .B1(output_p1_times_a1_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1712) );
  AOI32X1 U6275 ( .A0(n687), .A1(n1746), 
        .A2(output_p2_times_a2_div_componentxUDxcentral_parallel_output_0), 
        .B0(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[1]), 
        .B1(output_p2_times_a2_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1744) );
  OAI221XL U6276 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_8), 
        .A1(input_times_b0_div_componentxn53), 
        .B0(input_times_b0_div_componentxUDxcentral_parallel_output_9), 
        .B1(input_times_b0_div_componentxn54), .C0(n1546), .Y(n1547) );
  OAI221XL U6277 ( .A0(n853), .A1(n1531), .B0(n854), .B1(n1530), .C0(n1545), 
        .Y(n1546) );
  INVX1 U6278 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1530) );
  INVX1 U6279 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_7), 
        .Y(n1531) );
  OAI221XL U6280 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_8), 
        .A1(n4231), 
        .B0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_9), 
        .B1(n4232), .C0(n1622), .Y(n1623) );
  OAI221XL U6281 ( .A0(n1012), .A1(n1515), .B0(n1013), .B1(n1514), .C0(n1621), 
        .Y(n1622) );
  INVX1 U6282 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1514) );
  INVX1 U6283 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_7), 
        .Y(n1515) );
  OAI221XL U6284 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_8), 
        .A1(n4287), 
        .B0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_9), 
        .B1(n4288), .C0(n1603), .Y(n1604) );
  OAI221XL U6285 ( .A0(n1171), .A1(n1499), .B0(n1172), .B1(n1498), .C0(n1602), 
        .Y(n1603) );
  INVX1 U6286 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1498) );
  INVX1 U6287 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_7), 
        .Y(n1499) );
  OAI221XL U6288 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_8), 
        .A1(n4341), 
        .B0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_9), 
        .B1(n4342), .C0(n1584), .Y(n1585) );
  OAI221XL U6289 ( .A0(n535), .A1(n1483), .B0(n536), .B1(n1482), .C0(n1583), 
        .Y(n1584) );
  INVX1 U6290 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1482) );
  INVX1 U6291 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_7), 
        .Y(n1483) );
  OAI221XL U6292 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_8), 
        .A1(n4397), 
        .B0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_9), 
        .B1(n4398), .C0(n1565), .Y(n1566) );
  OAI221XL U6293 ( .A0(n694), .A1(n1467), .B0(n695), .B1(n1466), .C0(n1564), 
        .Y(n1565) );
  INVX1 U6294 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1466) );
  INVX1 U6295 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_7), 
        .Y(n1467) );
  OAI221XL U6296 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_2), 
        .A1(input_times_b0_div_componentxn47), 
        .B0(input_times_b0_div_componentxUDxcentral_parallel_output_3), 
        .B1(input_times_b0_div_componentxn48), .C0(n1540), .Y(n1541) );
  OAI222XL U6297 ( .A0(n1539), .A1(n1537), .B0(n847), .B1(n1538), .C0(n848), 
        .C1(n1536), .Y(n1540) );
  INVX1 U6298 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1536) );
  INVX1 U6299 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1537) );
  OAI221XL U6300 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_2), 
        .A1(n4225), 
        .B0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_3), 
        .B1(n4226), .C0(n1616), .Y(n1617) );
  OAI222XL U6301 ( .A0(n1615), .A1(n1521), .B0(n1006), .B1(n1614), .C0(n1007), 
        .C1(n1520), .Y(n1616) );
  INVX1 U6302 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1520) );
  INVX1 U6303 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1521) );
  OAI221XL U6304 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_2), 
        .A1(n4281), 
        .B0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_3), 
        .B1(n4282), .C0(n1597), .Y(n1598) );
  OAI222XL U6305 ( .A0(n1596), .A1(n1505), .B0(n1165), .B1(n1595), .C0(n1166), 
        .C1(n1504), .Y(n1597) );
  INVX1 U6306 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1504) );
  INVX1 U6307 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1505) );
  OAI221XL U6308 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_2), 
        .A1(n4335), 
        .B0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_3), 
        .B1(n4336), .C0(n1578), .Y(n1579) );
  OAI222XL U6309 ( .A0(n1577), .A1(n1489), .B0(n529), .B1(n1576), .C0(n530), 
        .C1(n1488), .Y(n1578) );
  INVX1 U6310 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1488) );
  INVX1 U6311 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1489) );
  OAI221XL U6312 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_2), 
        .A1(n4391), 
        .B0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_3), 
        .B1(n4392), .C0(n1559), .Y(n1560) );
  OAI222XL U6313 ( .A0(n1558), .A1(n1473), .B0(n688), .B1(n1557), .C0(n689), 
        .C1(n1472), .Y(n1559) );
  INVX1 U6314 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1472) );
  INVX1 U6315 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1473) );
  OAI221XL U6316 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_4), 
        .A1(input_times_b0_div_componentxn49), 
        .B0(input_times_b0_div_componentxUDxcentral_parallel_output_5), 
        .B1(input_times_b0_div_componentxn50), .C0(n1542), .Y(n1543) );
  OAI221XL U6317 ( .A0(n849), .A1(n1535), .B0(n850), .B1(n1534), .C0(n1541), 
        .Y(n1542) );
  INVX1 U6318 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1534) );
  INVX1 U6319 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_3), 
        .Y(n1535) );
  OAI221XL U6320 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_4), 
        .A1(n4227), 
        .B0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_5), 
        .B1(n4228), .C0(n1618), .Y(n1619) );
  OAI221XL U6321 ( .A0(n1008), .A1(n1519), .B0(n1009), .B1(n1518), .C0(n1617), 
        .Y(n1618) );
  INVX1 U6322 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1518) );
  INVX1 U6323 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_3), 
        .Y(n1519) );
  OAI221XL U6324 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_4), 
        .A1(n4283), 
        .B0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_5), 
        .B1(n4284), .C0(n1599), .Y(n1600) );
  OAI221XL U6325 ( .A0(n1167), .A1(n1503), .B0(n1168), .B1(n1502), .C0(n1598), 
        .Y(n1599) );
  INVX1 U6326 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1502) );
  INVX1 U6327 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_3), 
        .Y(n1503) );
  OAI221XL U6328 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_4), 
        .A1(n4337), 
        .B0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_5), 
        .B1(n4338), .C0(n1580), .Y(n1581) );
  OAI221XL U6329 ( .A0(n531), .A1(n1487), .B0(n532), .B1(n1486), .C0(n1579), 
        .Y(n1580) );
  INVX1 U6330 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1486) );
  INVX1 U6331 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_3), 
        .Y(n1487) );
  OAI221XL U6332 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_4), 
        .A1(n4393), 
        .B0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_5), 
        .B1(n4394), .C0(n1561), .Y(n1562) );
  OAI221XL U6333 ( .A0(n690), .A1(n1471), .B0(n691), .B1(n1470), .C0(n1560), 
        .Y(n1561) );
  INVX1 U6334 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1470) );
  INVX1 U6335 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_3), 
        .Y(n1471) );
  OAI221XL U6336 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_6), 
        .A1(input_times_b0_div_componentxn51), 
        .B0(input_times_b0_div_componentxUDxcentral_parallel_output_7), 
        .B1(input_times_b0_div_componentxn52), .C0(n1544), .Y(n1545) );
  OAI221XL U6337 ( .A0(n851), .A1(n1533), .B0(n852), .B1(n1532), .C0(n1543), 
        .Y(n1544) );
  INVX1 U6338 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1532) );
  INVX1 U6339 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_5), 
        .Y(n1533) );
  OAI221XL U6340 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_6), 
        .A1(n4229), 
        .B0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_7), 
        .B1(n4230), .C0(n1620), .Y(n1621) );
  OAI221XL U6341 ( .A0(n1010), .A1(n1517), .B0(n1011), .B1(n1516), .C0(n1619), 
        .Y(n1620) );
  INVX1 U6342 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1516) );
  INVX1 U6343 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_5), 
        .Y(n1517) );
  OAI221XL U6344 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_6), 
        .A1(n4285), 
        .B0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_7), 
        .B1(n4286), .C0(n1601), .Y(n1602) );
  OAI221XL U6345 ( .A0(n1169), .A1(n1501), .B0(n1170), .B1(n1500), .C0(n1600), 
        .Y(n1601) );
  INVX1 U6346 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1500) );
  INVX1 U6347 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_5), 
        .Y(n1501) );
  OAI221XL U6348 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_6), 
        .A1(n4339), 
        .B0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_7), 
        .B1(n4340), .C0(n1582), .Y(n1583) );
  OAI221XL U6349 ( .A0(n533), .A1(n1485), .B0(n534), .B1(n1484), .C0(n1581), 
        .Y(n1582) );
  INVX1 U6350 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1484) );
  INVX1 U6351 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_5), 
        .Y(n1485) );
  OAI221XL U6352 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_6), 
        .A1(n4395), 
        .B0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_7), 
        .B1(n4396), .C0(n1563), .Y(n1564) );
  OAI221XL U6353 ( .A0(n692), .A1(n1469), .B0(n693), .B1(n1468), .C0(n1562), 
        .Y(n1563) );
  INVX1 U6354 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1468) );
  INVX1 U6355 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_5), 
        .Y(n1469) );
  OAI221XL U6356 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_10), 
        .A1(input_times_b0_div_componentxn55), 
        .B0(input_times_b0_div_componentxUDxcentral_parallel_output_11), 
        .B1(input_times_b0_div_componentxn56), .C0(n1548), .Y(n1549) );
  OAI221XL U6357 ( .A0(n845), .A1(n1528), .B0(n855), .B1(n1529), .C0(n1547), 
        .Y(n1548) );
  INVX1 U6358 ( .A(input_times_b0_div_componentxn54), .Y(n855) );
  INVX1 U6359 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1528) );
  OAI221XL U6360 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_10), 
        .A1(n4233), 
        .B0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_11), 
        .B1(n4234), .C0(n1624), .Y(n1625) );
  OAI221XL U6361 ( .A0(n1004), .A1(n1512), .B0(n1014), .B1(n1513), .C0(n1623), 
        .Y(n1624) );
  INVX1 U6362 ( .A(n4232), .Y(n1014) );
  INVX1 U6363 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1512) );
  OAI221XL U6364 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_10), 
        .A1(n4289), 
        .B0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_11), 
        .B1(n4290), .C0(n1605), .Y(n1606) );
  OAI221XL U6365 ( .A0(n1163), .A1(n1496), .B0(n1173), .B1(n1497), .C0(n1604), 
        .Y(n1605) );
  INVX1 U6366 ( .A(n4288), .Y(n1173) );
  INVX1 U6367 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1496) );
  OAI221XL U6368 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_10), 
        .A1(n4343), 
        .B0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_11), 
        .B1(n4344), .C0(n1586), .Y(n1587) );
  OAI221XL U6369 ( .A0(n527), .A1(n1480), .B0(n537), .B1(n1481), .C0(n1585), 
        .Y(n1586) );
  INVX1 U6370 ( .A(n4342), .Y(n537) );
  INVX1 U6371 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1480) );
  OAI221XL U6372 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_10), 
        .A1(n4399), 
        .B0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_11), 
        .B1(n4400), .C0(n1567), .Y(n1568) );
  OAI221XL U6373 ( .A0(n686), .A1(n1464), .B0(n696), .B1(n1465), .C0(n1566), 
        .Y(n1567) );
  INVX1 U6374 ( .A(n4398), .Y(n696) );
  INVX1 U6375 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1464) );
  OAI221XL U6376 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_12), 
        .A1(input_times_b0_div_componentxn57), 
        .B0(input_times_b0_div_componentxUDxcentral_parallel_output_13), 
        .B1(input_times_b0_div_componentxn58), .C0(n1550), .Y(n1551) );
  OAI221XL U6377 ( .A0(n838), .A1(n1527), .B0(n839), .B1(n1526), .C0(n1549), 
        .Y(n1550) );
  INVX1 U6378 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1526) );
  INVX1 U6379 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_11), 
        .Y(n1527) );
  OAI221XL U6380 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_12), 
        .A1(n4235), 
        .B0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_13), 
        .B1(n4236), .C0(n1626), .Y(n1627) );
  OAI221XL U6381 ( .A0(n997), .A1(n1511), .B0(n998), .B1(n1510), .C0(n1625), 
        .Y(n1626) );
  INVX1 U6382 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1510) );
  INVX1 U6383 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_11), 
        .Y(n1511) );
  OAI221XL U6384 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_12), 
        .A1(n4291), 
        .B0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_13), 
        .B1(n4292), .C0(n1607), .Y(n1608) );
  OAI221XL U6385 ( .A0(n1156), .A1(n1495), .B0(n1157), .B1(n1494), .C0(n1606), 
        .Y(n1607) );
  INVX1 U6386 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1494) );
  INVX1 U6387 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_11), 
        .Y(n1495) );
  OAI221XL U6388 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_12), 
        .A1(n4345), 
        .B0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_13), 
        .B1(n4346), .C0(n1588), .Y(n1589) );
  OAI221XL U6389 ( .A0(n520), .A1(n1479), .B0(n521), .B1(n1478), .C0(n1587), 
        .Y(n1588) );
  INVX1 U6390 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1478) );
  INVX1 U6391 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_11), 
        .Y(n1479) );
  OAI221XL U6392 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_12), 
        .A1(n4401), 
        .B0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_13), 
        .B1(n4402), .C0(n1569), .Y(n1570) );
  OAI221XL U6393 ( .A0(n679), .A1(n1463), .B0(n680), .B1(n1462), .C0(n1568), 
        .Y(n1569) );
  INVX1 U6394 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1462) );
  INVX1 U6395 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_11), 
        .Y(n1463) );
  OAI221XL U6396 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_14), 
        .A1(input_times_b0_div_componentxn59), 
        .B0(input_times_b0_div_componentxUDxcentral_parallel_output_15), 
        .B1(input_times_b0_div_componentxn60), .C0(n1552), .Y(n1553) );
  OAI221XL U6397 ( .A0(n840), .A1(n1525), .B0(n841), .B1(n1524), .C0(n1551), 
        .Y(n1552) );
  INVX1 U6398 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1524) );
  INVX1 U6399 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_13), 
        .Y(n1525) );
  OAI221XL U6400 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_14), 
        .A1(n4237), 
        .B0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_15), 
        .B1(n4238), .C0(n1628), .Y(n1629) );
  OAI221XL U6401 ( .A0(n999), .A1(n1509), .B0(n1000), .B1(n1508), .C0(n1627), 
        .Y(n1628) );
  INVX1 U6402 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1508) );
  INVX1 U6403 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_13), 
        .Y(n1509) );
  OAI221XL U6404 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_14), 
        .A1(n4293), 
        .B0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_15), 
        .B1(n4294), .C0(n1609), .Y(n1610) );
  OAI221XL U6405 ( .A0(n1158), .A1(n1493), .B0(n1159), .B1(n1492), .C0(n1608), 
        .Y(n1609) );
  INVX1 U6406 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1492) );
  INVX1 U6407 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_13), 
        .Y(n1493) );
  OAI221XL U6408 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_14), 
        .A1(n4347), 
        .B0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_15), 
        .B1(n4348), .C0(n1590), .Y(n1591) );
  OAI221XL U6409 ( .A0(n522), .A1(n1477), .B0(n523), .B1(n1476), .C0(n1589), 
        .Y(n1590) );
  INVX1 U6410 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1476) );
  INVX1 U6411 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_13), 
        .Y(n1477) );
  OAI221XL U6412 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_14), 
        .A1(n4403), 
        .B0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_15), 
        .B1(n4404), .C0(n1571), .Y(n1572) );
  OAI221XL U6413 ( .A0(n681), .A1(n1461), .B0(n682), .B1(n1460), .C0(n1570), 
        .Y(n1571) );
  INVX1 U6414 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1460) );
  INVX1 U6415 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_13), 
        .Y(n1461) );
  AOI22X1 U6416 ( 
        .A0(input_times_b0_div_componentxUDxsub_ready_negative_divisor[3]), 
        .A1(input_times_b0_div_componentxUDxcentral_parallel_output_3), 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn13), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn14), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn12) );
  AOI22X1 U6417 ( 
        .A0(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[3]), 
        .A1(input_p1_times_b1_div_componentxUDxcentral_parallel_output_3), 
        .B0(n1645), .B1(n1646), .Y(n1644) );
  AOI22X1 U6418 ( 
        .A0(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[3]), 
        .A1(input_p2_times_b2_div_componentxUDxcentral_parallel_output_3), 
        .B0(n1677), .B1(n1678), .Y(n1676) );
  AOI22X1 U6419 ( 
        .A0(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[3]), 
        .A1(output_p1_times_a1_div_componentxUDxcentral_parallel_output_3), 
        .B0(n1709), .B1(n1710), .Y(n1708) );
  AOI22X1 U6420 ( 
        .A0(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[3]), 
        .A1(output_p2_times_a2_div_componentxUDxcentral_parallel_output_3), 
        .B0(n1741), .B1(n1742), .Y(n1740) );
  AOI22X1 U6421 ( 
        .A0(input_times_b0_div_componentxUDxsub_ready_negative_divisor[5]), 
        .A1(input_times_b0_div_componentxUDxcentral_parallel_output_5), 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn9), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn10), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn8) );
  AOI22X1 U6422 ( 
        .A0(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[5]), 
        .A1(input_p1_times_b1_div_componentxUDxcentral_parallel_output_5), 
        .B0(n1641), .B1(n1642), .Y(n1640) );
  AOI22X1 U6423 ( 
        .A0(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[5]), 
        .A1(input_p2_times_b2_div_componentxUDxcentral_parallel_output_5), 
        .B0(n1673), .B1(n1674), .Y(n1672) );
  AOI22X1 U6424 ( 
        .A0(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[5]), 
        .A1(output_p1_times_a1_div_componentxUDxcentral_parallel_output_5), 
        .B0(n1705), .B1(n1706), .Y(n1704) );
  AOI22X1 U6425 ( 
        .A0(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[5]), 
        .A1(output_p2_times_a2_div_componentxUDxcentral_parallel_output_5), 
        .B0(n1737), .B1(n1738), .Y(n1736) );
  AOI22X1 U6426 ( 
        .A0(input_times_b0_div_componentxUDxsub_ready_negative_divisor[7]), 
        .A1(input_times_b0_div_componentxUDxcentral_parallel_output_7), 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn5), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn6), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn4) );
  AOI22X1 U6427 ( 
        .A0(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[7]), 
        .A1(input_p1_times_b1_div_componentxUDxcentral_parallel_output_7), 
        .B0(n1637), .B1(n1638), .Y(n1636) );
  AOI22X1 U6428 ( 
        .A0(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[7]), 
        .A1(input_p2_times_b2_div_componentxUDxcentral_parallel_output_7), 
        .B0(n1669), .B1(n1670), .Y(n1668) );
  AOI22X1 U6429 ( 
        .A0(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[7]), 
        .A1(output_p1_times_a1_div_componentxUDxcentral_parallel_output_7), 
        .B0(n1701), .B1(n1702), .Y(n1700) );
  AOI22X1 U6430 ( 
        .A0(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[7]), 
        .A1(output_p2_times_a2_div_componentxUDxcentral_parallel_output_7), 
        .B0(n1733), .B1(n1734), .Y(n1732) );
  AOI22X1 U6431 ( 
        .A0(input_times_b0_div_componentxUDxsub_ready_negative_divisor[9]), 
        .A1(input_times_b0_div_componentxUDxcentral_parallel_output_9), 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn1), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn2), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn35) );
  AOI22X1 U6432 ( 
        .A0(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[9]), 
        .A1(input_p1_times_b1_div_componentxUDxcentral_parallel_output_9), 
        .B0(n1633), .B1(n1634), .Y(n1663) );
  AOI22X1 U6433 ( 
        .A0(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[9]), 
        .A1(input_p2_times_b2_div_componentxUDxcentral_parallel_output_9), 
        .B0(n1665), .B1(n1666), .Y(n1695) );
  AOI22X1 U6434 ( 
        .A0(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[9]), 
        .A1(output_p1_times_a1_div_componentxUDxcentral_parallel_output_9), 
        .B0(n1697), .B1(n1698), .Y(n1727) );
  AOI22X1 U6435 ( 
        .A0(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[9]), 
        .A1(output_p2_times_a2_div_componentxUDxcentral_parallel_output_9), 
        .B0(n1729), .B1(n1730), .Y(n1759) );
  AOI22X1 U6436 ( 
        .A0(input_times_b0_div_componentxUDxsub_ready_negative_divisor[11]), 
        .A1(input_times_b0_div_componentxUDxcentral_parallel_output_11), 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn33), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn34), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn31) );
  AOI22X1 U6437 ( 
        .A0(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[11]), 
        .A1(input_p1_times_b1_div_componentxUDxcentral_parallel_output_11), 
        .B0(n1661), .B1(n1662), .Y(n1659) );
  AOI22X1 U6438 ( 
        .A0(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[11]), 
        .A1(input_p2_times_b2_div_componentxUDxcentral_parallel_output_11), 
        .B0(n1693), .B1(n1694), .Y(n1691) );
  AOI22X1 U6439 ( 
        .A0(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[11]), 
        .A1(output_p1_times_a1_div_componentxUDxcentral_parallel_output_11), 
        .B0(n1725), .B1(n1726), .Y(n1723) );
  AOI22X1 U6440 ( 
        .A0(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[11]), 
        .A1(output_p2_times_a2_div_componentxUDxcentral_parallel_output_11), 
        .B0(n1757), .B1(n1758), .Y(n1755) );
  AOI22X1 U6441 ( 
        .A0(input_times_b0_div_componentxUDxsub_ready_negative_divisor[13]), 
        .A1(input_times_b0_div_componentxUDxcentral_parallel_output_13), 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn29), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn30), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn27) );
  AOI22X1 U6442 ( 
        .A0(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[13]), 
        .A1(input_p1_times_b1_div_componentxUDxcentral_parallel_output_13), 
        .B0(n1657), .B1(n1658), .Y(n1655) );
  AOI22X1 U6443 ( 
        .A0(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[13]), 
        .A1(input_p2_times_b2_div_componentxUDxcentral_parallel_output_13), 
        .B0(n1689), .B1(n1690), .Y(n1687) );
  AOI22X1 U6444 ( 
        .A0(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[13]), 
        .A1(output_p1_times_a1_div_componentxUDxcentral_parallel_output_13), 
        .B0(n1721), .B1(n1722), .Y(n1719) );
  AOI22X1 U6445 ( 
        .A0(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[13]), 
        .A1(output_p2_times_a2_div_componentxUDxcentral_parallel_output_13), 
        .B0(n1753), .B1(n1754), .Y(n1751) );
  OAI2BB2X1 U6446 ( 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn16), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn15), 
        .A0N(input_times_b0_div_componentxUDxsub_ready_negative_divisor[2]), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_2), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn13) );
  OAI2BB2X1 U6447 ( .B0(n1648), .B1(n1647), 
        .A0N(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[2]), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1645) );
  OAI2BB2X1 U6448 ( .B0(n1680), .B1(n1679), 
        .A0N(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[2]), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1677) );
  OAI2BB2X1 U6449 ( .B0(n1712), .B1(n1711), 
        .A0N(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[2]), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1709) );
  OAI2BB2X1 U6450 ( .B0(n1744), .B1(n1743), 
        .A0N(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[2]), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_2), 
        .Y(n1741) );
  OAI2BB2X1 U6451 ( 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn12), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn11), 
        .A0N(input_times_b0_div_componentxUDxsub_ready_negative_divisor[4]), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_4), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn9) );
  OAI2BB2X1 U6452 ( .B0(n1644), .B1(n1643), 
        .A0N(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[4]), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1641) );
  OAI2BB2X1 U6453 ( .B0(n1676), .B1(n1675), 
        .A0N(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[4]), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1673) );
  OAI2BB2X1 U6454 ( .B0(n1708), .B1(n1707), 
        .A0N(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[4]), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1705) );
  OAI2BB2X1 U6455 ( .B0(n1740), .B1(n1739), 
        .A0N(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[4]), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_4), 
        .Y(n1737) );
  OAI2BB2X1 U6456 ( 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn8), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn7), 
        .A0N(input_times_b0_div_componentxUDxsub_ready_negative_divisor[6]), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_6), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn5) );
  OAI2BB2X1 U6457 ( .B0(n1640), .B1(n1639), 
        .A0N(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[6]), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1637) );
  OAI2BB2X1 U6458 ( .B0(n1672), .B1(n1671), 
        .A0N(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[6]), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1669) );
  OAI2BB2X1 U6459 ( .B0(n1704), .B1(n1703), 
        .A0N(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[6]), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1701) );
  OAI2BB2X1 U6460 ( .B0(n1736), .B1(n1735), 
        .A0N(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[6]), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_6), 
        .Y(n1733) );
  OAI2BB2X1 U6461 ( 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn4), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn3), 
        .A0N(input_times_b0_div_componentxUDxsub_ready_negative_divisor[8]), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_8), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn1) );
  OAI2BB2X1 U6462 ( .B0(n1636), .B1(n1635), 
        .A0N(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[8]), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1633) );
  OAI2BB2X1 U6463 ( .B0(n1668), .B1(n1667), 
        .A0N(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[8]), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1665) );
  OAI2BB2X1 U6464 ( .B0(n1700), .B1(n1699), 
        .A0N(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[8]), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1697) );
  OAI2BB2X1 U6465 ( .B0(n1732), .B1(n1731), 
        .A0N(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[8]), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_8), 
        .Y(n1729) );
  OAI2BB2X1 U6466 ( 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn35), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn36), 
        .A0N(input_times_b0_div_componentxUDxsub_ready_negative_divisor[10]), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_10), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn33) );
  OAI2BB2X1 U6467 ( .B0(n1663), .B1(n1664), 
        .A0N(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[10]), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1661) );
  OAI2BB2X1 U6468 ( .B0(n1695), .B1(n1696), 
        .A0N(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[10]), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1693) );
  OAI2BB2X1 U6469 ( .B0(n1727), .B1(n1728), 
        .A0N(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[10]), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1725) );
  OAI2BB2X1 U6470 ( .B0(n1759), .B1(n1760), 
        .A0N(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[10]), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_10), 
        .Y(n1757) );
  OAI2BB2X1 U6471 ( 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn31), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn32), 
        .A0N(input_times_b0_div_componentxUDxsub_ready_negative_divisor[12]), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_12), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn29) );
  OAI2BB2X1 U6472 ( .B0(n1659), .B1(n1660), 
        .A0N(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[12]), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1657) );
  OAI2BB2X1 U6473 ( .B0(n1691), .B1(n1692), 
        .A0N(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[12]), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1689) );
  OAI2BB2X1 U6474 ( .B0(n1723), .B1(n1724), 
        .A0N(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[12]), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1721) );
  OAI2BB2X1 U6475 ( .B0(n1755), .B1(n1756), 
        .A0N(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[12]), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_12), 
        .Y(n1753) );
  OAI2BB2X1 U6476 ( 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn27), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn28), 
        .A0N(input_times_b0_div_componentxUDxsub_ready_negative_divisor[14]), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_14), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn25) );
  OAI2BB2X1 U6477 ( .B0(n1655), .B1(n1656), 
        .A0N(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[14]), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1653) );
  OAI2BB2X1 U6478 ( .B0(n1687), .B1(n1688), 
        .A0N(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[14]), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1685) );
  OAI2BB2X1 U6479 ( .B0(n1719), .B1(n1720), 
        .A0N(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[14]), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1717) );
  OAI2BB2X1 U6480 ( .B0(n1751), .B1(n1752), 
        .A0N(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[14]), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_14), 
        .Y(n1749) );
  AOI22X1 U6481 ( 
        .A0(input_times_b0_div_componentxUDxsub_ready_negative_divisor[15]), 
        .A1(input_times_b0_div_componentxUDxcentral_parallel_output_15), 
        .B0(input_times_b0_div_componentxUDxactually_substractsxn25), 
        .B1(input_times_b0_div_componentxUDxactually_substractsxn26), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn23) );
  AOI22X1 U6482 ( 
        .A0(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[15]), 
        .A1(input_p1_times_b1_div_componentxUDxcentral_parallel_output_15), 
        .B0(n1653), .B1(n1654), .Y(n1651) );
  AOI22X1 U6483 ( 
        .A0(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[15]), 
        .A1(input_p2_times_b2_div_componentxUDxcentral_parallel_output_15), 
        .B0(n1685), .B1(n1686), .Y(n1683) );
  AOI22X1 U6484 ( 
        .A0(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[15]), 
        .A1(output_p1_times_a1_div_componentxUDxcentral_parallel_output_15), 
        .B0(n1717), .B1(n1718), .Y(n1715) );
  AOI22X1 U6485 ( 
        .A0(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[15]), 
        .A1(output_p2_times_a2_div_componentxUDxcentral_parallel_output_15), 
        .B0(n1749), .B1(n1750), .Y(n1747) );
  XOR2X1 U6486 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_3), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[3]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn14) );
  XOR2X1 U6487 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_3), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[3]), 
        .Y(n1646) );
  XOR2X1 U6488 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_3), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[3]), 
        .Y(n1678) );
  XOR2X1 U6489 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_3), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[3]), 
        .Y(n1710) );
  XOR2X1 U6490 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_3), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[3]), 
        .Y(n1742) );
  NOR2BX1 U6491 ( .AN(n846), 
        .B(input_times_b0_div_componentxUDxcentral_parallel_output_0), 
        .Y(n1539) );
  NOR2BX1 U6492 ( .AN(n1005), 
        .B(input_p1_times_b1_div_componentxUDxcentral_parallel_output_0), 
        .Y(n1615) );
  NOR2BX1 U6493 ( .AN(n1164), 
        .B(input_p2_times_b2_div_componentxUDxcentral_parallel_output_0), 
        .Y(n1596) );
  NOR2BX1 U6494 ( .AN(n528), 
        .B(output_p1_times_a1_div_componentxUDxcentral_parallel_output_0), 
        .Y(n1577) );
  NOR2BX1 U6495 ( .AN(n687), 
        .B(output_p2_times_a2_div_componentxUDxcentral_parallel_output_0), 
        .Y(n1558) );
  OAI2BB2X1 U6496 ( .B0(n1236), .B1(n1260), 
        .A0N(output_p2_times_a2_mul_componentxinput_A_inverted[0]), .A1N(n320), 
        .Y(n4655) );
  INVX1 U6497 ( .A(\output_signal[0] ), .Y(n1236) );
  OAI2BB2X1 U6498 ( .B0(n1226), .B1(n1260), .A0N(output_previous_2[1]), 
        .A1N(n320), .Y(n4656) );
  XOR2X1 U6499 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_1), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[1]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn18) );
  XOR2X1 U6500 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_1), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[1]), 
        .Y(n1650) );
  XOR2X1 U6501 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_1), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[1]), 
        .Y(n1682) );
  XOR2X1 U6502 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_1), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[1]), 
        .Y(n1714) );
  XOR2X1 U6503 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_1), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[1]), 
        .Y(n1746) );
  XNOR2X1 U6504 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_2), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[2]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn15) );
  XNOR2X1 U6505 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_2), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[2]), 
        .Y(n1647) );
  XNOR2X1 U6506 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_2), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[2]), 
        .Y(n1679) );
  XNOR2X1 U6507 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_2), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[2]), 
        .Y(n1711) );
  XNOR2X1 U6508 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_2), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[2]), 
        .Y(n1743) );
  OAI2BB2X1 U6509 ( .B0(n1212), .B1(n320), .A0N(output_previous_2[8]), 
        .A1N(n320), .Y(n4663) );
  INVX1 U6510 ( .A(output_previous_1[8]), .Y(n1212) );
  NOR2BX1 U6511 ( .AN(n1539), 
        .B(input_times_b0_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1538) );
  NOR2BX1 U6512 ( .AN(n1615), 
        .B(input_p1_times_b1_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1614) );
  NOR2BX1 U6513 ( .AN(n1596), 
        .B(input_p2_times_b2_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1595) );
  NOR2BX1 U6514 ( .AN(n1577), 
        .B(output_p1_times_a1_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1576) );
  NOR2BX1 U6515 ( .AN(n1558), 
        .B(output_p2_times_a2_div_componentxUDxcentral_parallel_output_1), 
        .Y(n1557) );
  OAI2BB1X1 U6516 ( .A0N(n1522), .A1N(n843), .B0(n1554), .Y(n1555) );
  OAI221XL U6517 ( .A0(n842), .A1(n1523), .B0(n843), .B1(n1522), .C0(n1553), 
        .Y(n1554) );
  INVX1 U6518 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_16), 
        .Y(n1522) );
  INVX1 U6519 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_15), 
        .Y(n1523) );
  OAI2BB1X1 U6520 ( .A0N(n1506), .A1N(n1002), .B0(n1630), .Y(n1631) );
  OAI221XL U6521 ( .A0(n1001), .A1(n1507), .B0(n1002), .B1(n1506), .C0(n1629), 
        .Y(n1630) );
  INVX1 U6522 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_16), 
        .Y(n1506) );
  INVX1 U6523 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_15), 
        .Y(n1507) );
  OAI2BB1X1 U6524 ( .A0N(n1490), .A1N(n1161), .B0(n1611), .Y(n1612) );
  OAI221XL U6525 ( .A0(n1160), .A1(n1491), .B0(n1161), .B1(n1490), .C0(n1610), 
        .Y(n1611) );
  INVX1 U6526 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_16), 
        .Y(n1490) );
  INVX1 U6527 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_15), 
        .Y(n1491) );
  OAI2BB1X1 U6528 ( .A0N(n1474), .A1N(n525), .B0(n1592), .Y(n1593) );
  OAI221XL U6529 ( .A0(n524), .A1(n1475), .B0(n525), .B1(n1474), .C0(n1591), 
        .Y(n1592) );
  INVX1 U6530 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_16), 
        .Y(n1474) );
  INVX1 U6531 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_15), 
        .Y(n1475) );
  OAI2BB1X1 U6532 ( .A0N(n1458), .A1N(n684), .B0(n1573), .Y(n1574) );
  OAI221XL U6533 ( .A0(n683), .A1(n1459), .B0(n684), .B1(n1458), .C0(n1572), 
        .Y(n1573) );
  INVX1 U6534 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_16), 
        .Y(n1458) );
  INVX1 U6535 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_15), 
        .Y(n1459) );
  INVX1 U6536 ( .A(input_times_b0_div_componentxUDxis_less_than), .Y(n837) );
  OAI21XL U6537 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_17), 
        .A1(n844), .B0(n1556), 
        .Y(input_times_b0_div_componentxUDxis_less_than) );
  OAI2BB1X1 U6538 ( .A0N(n844), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_17), 
        .B0(n1555), .Y(n1556) );
  INVX1 U6539 ( .A(input_times_b0_div_componentxunsigned_B_17), .Y(n844) );
  INVX1 U6540 ( .A(input_p1_times_b1_div_componentxUDxis_less_than), .Y(n996)
         );
  OAI21XL U6541 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_17), 
        .A1(n1003), .B0(n1632), 
        .Y(input_p1_times_b1_div_componentxUDxis_less_than) );
  OAI2BB1X1 U6542 ( .A0N(n1003), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_17), 
        .B0(n1631), .Y(n1632) );
  INVX1 U6543 ( .A(input_p1_times_b1_div_componentxunsigned_B_17), .Y(n1003)
         );
  INVX1 U6544 ( .A(input_p2_times_b2_div_componentxUDxis_less_than), .Y(n1155)
         );
  OAI21XL U6545 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_17), 
        .A1(n1162), .B0(n1613), 
        .Y(input_p2_times_b2_div_componentxUDxis_less_than) );
  OAI2BB1X1 U6546 ( .A0N(n1162), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_17), 
        .B0(n1612), .Y(n1613) );
  INVX1 U6547 ( .A(input_p2_times_b2_div_componentxunsigned_B_17), .Y(n1162)
         );
  INVX1 U6548 ( .A(output_p1_times_a1_div_componentxUDxis_less_than), .Y(n519)
         );
  OAI21XL U6549 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_17), 
        .A1(n526), .B0(n1594), 
        .Y(output_p1_times_a1_div_componentxUDxis_less_than) );
  OAI2BB1X1 U6550 ( .A0N(n526), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_17), 
        .B0(n1593), .Y(n1594) );
  INVX1 U6551 ( .A(output_p1_times_a1_div_componentxunsigned_B_17), .Y(n526)
         );
  INVX1 U6552 ( .A(output_p2_times_a2_div_componentxUDxis_less_than), .Y(n678)
         );
  OAI21XL U6553 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_17), 
        .A1(n685), .B0(n1575), 
        .Y(output_p2_times_a2_div_componentxUDxis_less_than) );
  OAI2BB1X1 U6554 ( .A0N(n685), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_17), 
        .B0(n1574), .Y(n1575) );
  INVX1 U6555 ( .A(output_p2_times_a2_div_componentxunsigned_B_17), .Y(n685)
         );
  OAI2BB1X1 U6556 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_4), 
        .B0(n1810), .Y(n1828) );
  AOI22X1 U6557 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_3), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[3]), 
        .B1(n14), .Y(n1810) );
  XOR2X1 U6558 ( .A(input_times_b0_div_componentxUDxactually_substractsxn13), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn14), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[3]) );
  OAI2BB1X1 U6559 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_6), 
        .B0(n1808), .Y(n1826) );
  AOI22X1 U6560 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_5), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[5]), 
        .B1(n14), .Y(n1808) );
  XOR2X1 U6561 ( .A(input_times_b0_div_componentxUDxactually_substractsxn9), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn10), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[5]) );
  OAI2BB1X1 U6562 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_8), 
        .B0(n1806), .Y(n1824) );
  AOI22X1 U6563 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_7), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[7]), 
        .B1(n14), .Y(n1806) );
  XOR2X1 U6564 ( .A(input_times_b0_div_componentxUDxactually_substractsxn5), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn6), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[7]) );
  OAI2BB1X1 U6565 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_10), 
        .B0(n1804), .Y(n1822) );
  AOI22X1 U6566 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_9), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[9]), 
        .B1(n14), .Y(n1804) );
  XOR2X1 U6567 ( .A(input_times_b0_div_componentxUDxactually_substractsxn1), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn2), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[9]) );
  OAI2BB1X1 U6568 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_12), 
        .B0(n1802), .Y(n1820) );
  AOI22X1 U6569 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_11), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[11]), 
        .B1(n14), .Y(n1802) );
  XOR2X1 U6570 ( .A(input_times_b0_div_componentxUDxactually_substractsxn33), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn34), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[11])
         );
  OAI2BB1X1 U6571 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_14), 
        .B0(n1800), .Y(n1818) );
  AOI22X1 U6572 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_13), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[13]), 
        .B1(n14), .Y(n1800) );
  XOR2X1 U6573 ( .A(input_times_b0_div_componentxUDxactually_substractsxn29), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn30), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[13])
         );
  OAI2BB1X1 U6574 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_16), 
        .B0(n1798), .Y(n1816) );
  AOI22X1 U6575 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_15), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[15]), 
        .B1(n14), .Y(n1798) );
  XOR2X1 U6576 ( .A(input_times_b0_div_componentxUDxactually_substractsxn25), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn26), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[15])
         );
  OAI2BB1X1 U6577 ( .A0N(n367), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_4), 
        .B0(n1920), .Y(n1938) );
  AOI22X1 U6578 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_3), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[3]), 
        .B1(n15), .Y(n1920) );
  XOR2X1 U6579 ( .A(n1645), .B(n1646), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[3])
         );
  OAI2BB1X1 U6580 ( .A0N(n371), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_6), 
        .B0(n1918), .Y(n1936) );
  AOI22X1 U6581 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_5), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[5]), 
        .B1(n15), .Y(n1918) );
  XOR2X1 U6582 ( .A(n1641), .B(n1642), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[5])
         );
  OAI2BB1X1 U6583 ( .A0N(n368), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_8), 
        .B0(n1916), .Y(n1934) );
  AOI22X1 U6584 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_7), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[7]), 
        .B1(n15), .Y(n1916) );
  XOR2X1 U6585 ( .A(n1637), .B(n1638), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[7])
         );
  OAI2BB1X1 U6586 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_10), 
        .B0(n1914), .Y(n1932) );
  AOI22X1 U6587 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_9), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[9]), 
        .B1(n15), .Y(n1914) );
  XOR2X1 U6588 ( .A(n1633), .B(n1634), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[9])
         );
  OAI2BB1X1 U6589 ( .A0N(n372), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_12), 
        .B0(n1912), .Y(n1930) );
  AOI22X1 U6590 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_11), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[11]), 
        .B1(n15), .Y(n1912) );
  XOR2X1 U6591 ( .A(n1661), .B(n1662), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[11])
         );
  OAI2BB1X1 U6592 ( .A0N(n367), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_14), 
        .B0(n1910), .Y(n1928) );
  AOI22X1 U6593 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_13), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[13]), 
        .B1(n15), .Y(n1910) );
  XOR2X1 U6594 ( .A(n1657), .B(n1658), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[13])
         );
  OAI2BB1X1 U6595 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_16), 
        .B0(n1908), .Y(n1926) );
  AOI22X1 U6596 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_15), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[15]), 
        .B1(n15), .Y(n1908) );
  XOR2X1 U6597 ( .A(n1653), .B(n1654), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[15])
         );
  OAI2BB1X1 U6598 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_4), 
        .B0(n2029), .Y(n2047) );
  AOI22X1 U6599 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_3), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[3]), 
        .B1(n16), .Y(n2029) );
  XOR2X1 U6600 ( .A(n1677), .B(n1678), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[3])
         );
  OAI2BB1X1 U6601 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_6), 
        .B0(n2027), .Y(n2045) );
  AOI22X1 U6602 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_5), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[5]), 
        .B1(n16), .Y(n2027) );
  XOR2X1 U6603 ( .A(n1673), .B(n1674), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[5])
         );
  OAI2BB1X1 U6604 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_8), 
        .B0(n2025), .Y(n2043) );
  AOI22X1 U6605 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_7), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[7]), 
        .B1(n16), .Y(n2025) );
  XOR2X1 U6606 ( .A(n1669), .B(n1670), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[7])
         );
  OAI2BB1X1 U6607 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_10), 
        .B0(n2023), .Y(n2041) );
  AOI22X1 U6608 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_9), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[9]), 
        .B1(n16), .Y(n2023) );
  XOR2X1 U6609 ( .A(n1665), .B(n1666), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[9])
         );
  OAI2BB1X1 U6610 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_12), 
        .B0(n2021), .Y(n2039) );
  AOI22X1 U6611 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_11), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[11]), 
        .B1(n16), .Y(n2021) );
  XOR2X1 U6612 ( .A(n1693), .B(n1694), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[11])
         );
  OAI2BB1X1 U6613 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_14), 
        .B0(n2019), .Y(n2037) );
  AOI22X1 U6614 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_13), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[13]), 
        .B1(n16), .Y(n2019) );
  XOR2X1 U6615 ( .A(n1689), .B(n1690), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[13])
         );
  OAI2BB1X1 U6616 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_16), 
        .B0(n2017), .Y(n2035) );
  AOI22X1 U6617 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_15), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[15]), 
        .B1(n16), .Y(n2017) );
  XOR2X1 U6618 ( .A(n1685), .B(n1686), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[15])
         );
  OAI2BB1X1 U6619 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_4), 
        .B0(n2139), .Y(n2157) );
  AOI22X1 U6620 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_3), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[3]), 
        .B1(n17), .Y(n2139) );
  XOR2X1 U6621 ( .A(n1709), .B(n1710), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[3])
         );
  OAI2BB1X1 U6622 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_6), 
        .B0(n2137), .Y(n2155) );
  AOI22X1 U6623 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_5), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[5]), 
        .B1(n17), .Y(n2137) );
  XOR2X1 U6624 ( .A(n1705), .B(n1706), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[5])
         );
  OAI2BB1X1 U6625 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_8), 
        .B0(n2135), .Y(n2153) );
  AOI22X1 U6626 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_7), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[7]), 
        .B1(n17), .Y(n2135) );
  XOR2X1 U6627 ( .A(n1701), .B(n1702), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[7])
         );
  OAI2BB1X1 U6628 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_10), 
        .B0(n2133), .Y(n2151) );
  AOI22X1 U6629 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_9), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[9]), 
        .B1(n17), .Y(n2133) );
  XOR2X1 U6630 ( .A(n1697), .B(n1698), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[9])
         );
  OAI2BB1X1 U6631 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_12), 
        .B0(n2131), .Y(n2149) );
  AOI22X1 U6632 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_11), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[11]), 
        .B1(n17), .Y(n2131) );
  XOR2X1 U6633 ( .A(n1725), .B(n1726), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[11])
         );
  OAI2BB1X1 U6634 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_14), 
        .B0(n2129), .Y(n2147) );
  AOI22X1 U6635 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_13), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[13]), 
        .B1(n17), .Y(n2129) );
  XOR2X1 U6636 ( .A(n1721), .B(n1722), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[13])
         );
  OAI2BB1X1 U6637 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_16), 
        .B0(n2127), .Y(n2145) );
  AOI22X1 U6638 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_15), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[15]), 
        .B1(n17), .Y(n2127) );
  XOR2X1 U6639 ( .A(n1717), .B(n1718), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[15])
         );
  OAI2BB1X1 U6640 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_4), 
        .B0(n2248), .Y(n2266) );
  AOI22X1 U6641 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_3), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[3]), 
        .B1(n18), .Y(n2248) );
  XOR2X1 U6642 ( .A(n1741), .B(n1742), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[3])
         );
  OAI2BB1X1 U6643 ( .A0N(n368), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_6), 
        .B0(n2246), .Y(n2264) );
  AOI22X1 U6644 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_5), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[5]), 
        .B1(n18), .Y(n2246) );
  XOR2X1 U6645 ( .A(n1737), .B(n1738), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[5])
         );
  OAI2BB1X1 U6646 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_8), 
        .B0(n2244), .Y(n2262) );
  AOI22X1 U6647 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_7), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[7]), 
        .B1(n18), .Y(n2244) );
  XOR2X1 U6648 ( .A(n1733), .B(n1734), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[7])
         );
  OAI2BB1X1 U6649 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_10), 
        .B0(n2242), .Y(n2260) );
  AOI22X1 U6650 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_9), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[9]), 
        .B1(n18), .Y(n2242) );
  XOR2X1 U6651 ( .A(n1729), .B(n1730), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[9])
         );
  OAI2BB1X1 U6652 ( .A0N(n370), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_12), 
        .B0(n2240), .Y(n2258) );
  AOI22X1 U6653 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_11), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[11]), 
        .B1(n18), .Y(n2240) );
  XOR2X1 U6654 ( .A(n1757), .B(n1758), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[11])
         );
  OAI2BB1X1 U6655 ( .A0N(n369), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_14), 
        .B0(n2238), .Y(n2256) );
  AOI22X1 U6656 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_13), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[13]), 
        .B1(n18), .Y(n2238) );
  XOR2X1 U6657 ( .A(n1753), .B(n1754), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[13])
         );
  OAI2BB1X1 U6658 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_16), 
        .B0(n2236), .Y(n2254) );
  AOI22X1 U6659 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_15), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[15]), 
        .B1(n18), .Y(n2236) );
  XOR2X1 U6660 ( .A(n1749), .B(n1750), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[15])
         );
  OAI2BB1X1 U6661 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_2), 
        .B0(n1812), .Y(n1830) );
  AOI22X1 U6662 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_1), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[1]), 
        .B1(n14), .Y(n1812) );
  XOR2X1 U6663 ( .A(input_times_b0_div_componentxUDxactually_substractsxn17), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn18), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[1]) );
  AND2X2 U6664 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_0), 
        .B(n846), .Y(input_times_b0_div_componentxUDxactually_substractsxn17)
         );
  OAI2BB1X1 U6665 ( .A0N(n367), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_2), 
        .B0(n1922), .Y(n1940) );
  AOI22X1 U6666 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_1), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[1]), 
        .B1(n15), .Y(n1922) );
  XOR2X1 U6667 ( .A(n1649), .B(n1650), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[1])
         );
  AND2X2 U6668 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_0), 
        .B(n1005), .Y(n1649) );
  OAI2BB1X1 U6669 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_2), 
        .B0(n2031), .Y(n2049) );
  AOI22X1 U6670 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_1), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[1]), 
        .B1(n16), .Y(n2031) );
  XOR2X1 U6671 ( .A(n1681), .B(n1682), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[1])
         );
  AND2X2 U6672 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_0), 
        .B(n1164), .Y(n1681) );
  OAI2BB1X1 U6673 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_2), 
        .B0(n2141), .Y(n2159) );
  AOI22X1 U6674 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_1), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[1]), 
        .B1(n17), .Y(n2141) );
  XOR2X1 U6675 ( .A(n1713), .B(n1714), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[1])
         );
  AND2X2 U6676 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_0), 
        .B(n528), .Y(n1713) );
  OAI2BB1X1 U6677 ( .A0N(n367), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_2), 
        .B0(n2250), .Y(n2268) );
  AOI22X1 U6678 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_1), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[1]), 
        .B1(n18), .Y(n2250) );
  XOR2X1 U6679 ( .A(n1745), .B(n1746), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[1])
         );
  AND2X2 U6680 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_0), 
        .B(n687), .Y(n1745) );
  OAI2BB1X1 U6681 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_1), 
        .B0(n1813), .Y(n1831) );
  AOI22X1 U6682 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_0), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[0]), 
        .B1(n14), .Y(n1813) );
  XOR2X1 U6683 ( .A(n846), 
        .B(input_times_b0_div_componentxUDxcentral_parallel_output_0), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[0]) );
  OAI2BB1X1 U6684 ( .A0N(n371), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_1), 
        .B0(n1923), .Y(n1941) );
  AOI22X1 U6685 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_0), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[0]), 
        .B1(n15), .Y(n1923) );
  XOR2X1 U6686 ( .A(n1005), 
        .B(input_p1_times_b1_div_componentxUDxcentral_parallel_output_0), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[0])
         );
  OAI2BB1X1 U6687 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_1), 
        .B0(n2032), .Y(n2050) );
  AOI22X1 U6688 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_0), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[0]), 
        .B1(n16), .Y(n2032) );
  XOR2X1 U6689 ( .A(n1164), 
        .B(input_p2_times_b2_div_componentxUDxcentral_parallel_output_0), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[0])
         );
  OAI2BB1X1 U6690 ( .A0N(n367), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_1), 
        .B0(n2142), .Y(n2160) );
  AOI22X1 U6691 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_0), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[0]), 
        .B1(n17), .Y(n2142) );
  XOR2X1 U6692 ( .A(n528), 
        .B(output_p1_times_a1_div_componentxUDxcentral_parallel_output_0), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[0])
         );
  OAI2BB1X1 U6693 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_1), 
        .B0(n2251), .Y(n2269) );
  AOI22X1 U6694 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_0), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[0]), 
        .B1(n18), .Y(n2251) );
  XOR2X1 U6695 ( .A(n687), 
        .B(output_p2_times_a2_div_componentxUDxcentral_parallel_output_0), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[0])
         );
  OAI2BB1X1 U6696 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_3), 
        .B0(n1811), .Y(n1829) );
  AOI22X1 U6697 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_2), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[2]), 
        .B1(n14), .Y(n1811) );
  XOR2X1 U6698 ( .A(input_times_b0_div_componentxUDxactually_substractsxn15), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn16), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[2]) );
  OAI2BB1X1 U6699 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_5), 
        .B0(n1809), .Y(n1827) );
  AOI22X1 U6700 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_4), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[4]), 
        .B1(n14), .Y(n1809) );
  XOR2X1 U6701 ( .A(input_times_b0_div_componentxUDxactually_substractsxn11), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn12), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[4]) );
  OAI2BB1X1 U6702 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_7), 
        .B0(n1807), .Y(n1825) );
  AOI22X1 U6703 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_6), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[6]), 
        .B1(n14), .Y(n1807) );
  XOR2X1 U6704 ( .A(input_times_b0_div_componentxUDxactually_substractsxn7), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn8), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[6]) );
  OAI2BB1X1 U6705 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_9), 
        .B0(n1805), .Y(n1823) );
  AOI22X1 U6706 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_8), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[8]), 
        .B1(n14), .Y(n1805) );
  XOR2X1 U6707 ( .A(input_times_b0_div_componentxUDxactually_substractsxn3), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn4), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[8]) );
  OAI2BB1X1 U6708 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_11), 
        .B0(n1803), .Y(n1821) );
  AOI22X1 U6709 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_10), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[10]), 
        .B1(n14), .Y(n1803) );
  XOR2X1 U6710 ( .A(input_times_b0_div_componentxUDxactually_substractsxn36), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn35), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[10])
         );
  OAI2BB1X1 U6711 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_13), 
        .B0(n1801), .Y(n1819) );
  AOI22X1 U6712 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_12), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[12]), 
        .B1(n14), .Y(n1801) );
  XOR2X1 U6713 ( .A(input_times_b0_div_componentxUDxactually_substractsxn32), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn31), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[12])
         );
  OAI2BB1X1 U6714 ( .A0N(n371), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_15), 
        .B0(n1799), .Y(n1817) );
  AOI22X1 U6715 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_14), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[14]), 
        .B1(n14), .Y(n1799) );
  XOR2X1 U6716 ( .A(input_times_b0_div_componentxUDxactually_substractsxn28), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn27), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[14])
         );
  OAI2BB1X1 U6717 ( .A0N(n368), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_3), 
        .B0(n1921), .Y(n1939) );
  AOI22X1 U6718 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_2), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[2]), 
        .B1(n15), .Y(n1921) );
  XOR2X1 U6719 ( .A(n1647), .B(n1648), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[2])
         );
  OAI2BB1X1 U6720 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_5), 
        .B0(n1919), .Y(n1937) );
  AOI22X1 U6721 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_4), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[4]), 
        .B1(n15), .Y(n1919) );
  XOR2X1 U6722 ( .A(n1643), .B(n1644), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[4])
         );
  OAI2BB1X1 U6723 ( .A0N(n372), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_7), 
        .B0(n1917), .Y(n1935) );
  AOI22X1 U6724 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_6), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[6]), 
        .B1(n15), .Y(n1917) );
  XOR2X1 U6725 ( .A(n1639), .B(n1640), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[6])
         );
  OAI2BB1X1 U6726 ( .A0N(n368), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_9), 
        .B0(n1915), .Y(n1933) );
  AOI22X1 U6727 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_8), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[8]), 
        .B1(n15), .Y(n1915) );
  XOR2X1 U6728 ( .A(n1635), .B(n1636), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[8])
         );
  OAI2BB1X1 U6729 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_11), 
        .B0(n1913), .Y(n1931) );
  AOI22X1 U6730 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_10), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[10]), 
        .B1(n15), .Y(n1913) );
  XOR2X1 U6731 ( .A(n1664), .B(n1663), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[10])
         );
  OAI2BB1X1 U6732 ( .A0N(n367), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_13), 
        .B0(n1911), .Y(n1929) );
  AOI22X1 U6733 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_12), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[12]), 
        .B1(n15), .Y(n1911) );
  XOR2X1 U6734 ( .A(n1660), .B(n1659), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[12])
         );
  OAI2BB1X1 U6735 ( .A0N(n371), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_15), 
        .B0(n1909), .Y(n1927) );
  AOI22X1 U6736 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_14), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[14]), 
        .B1(n15), .Y(n1909) );
  XOR2X1 U6737 ( .A(n1656), .B(n1655), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[14])
         );
  OAI2BB1X1 U6738 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_3), 
        .B0(n2030), .Y(n2048) );
  AOI22X1 U6739 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_2), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[2]), 
        .B1(n16), .Y(n2030) );
  XOR2X1 U6740 ( .A(n1679), .B(n1680), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[2])
         );
  OAI2BB1X1 U6741 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_5), 
        .B0(n2028), .Y(n2046) );
  AOI22X1 U6742 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_4), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[4]), 
        .B1(n16), .Y(n2028) );
  XOR2X1 U6743 ( .A(n1675), .B(n1676), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[4])
         );
  OAI2BB1X1 U6744 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_7), 
        .B0(n2026), .Y(n2044) );
  AOI22X1 U6745 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_6), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[6]), 
        .B1(n16), .Y(n2026) );
  XOR2X1 U6746 ( .A(n1671), .B(n1672), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[6])
         );
  OAI2BB1X1 U6747 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_9), 
        .B0(n2024), .Y(n2042) );
  AOI22X1 U6748 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_8), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[8]), 
        .B1(n16), .Y(n2024) );
  XOR2X1 U6749 ( .A(n1667), .B(n1668), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[8])
         );
  OAI2BB1X1 U6750 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_11), 
        .B0(n2022), .Y(n2040) );
  AOI22X1 U6751 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_10), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[10]), 
        .B1(n16), .Y(n2022) );
  XOR2X1 U6752 ( .A(n1696), .B(n1695), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[10])
         );
  OAI2BB1X1 U6753 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_13), 
        .B0(n2020), .Y(n2038) );
  AOI22X1 U6754 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_12), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[12]), 
        .B1(n16), .Y(n2020) );
  XOR2X1 U6755 ( .A(n1692), .B(n1691), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[12])
         );
  OAI2BB1X1 U6756 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_15), 
        .B0(n2018), .Y(n2036) );
  AOI22X1 U6757 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_14), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[14]), 
        .B1(n16), .Y(n2018) );
  XOR2X1 U6758 ( .A(n1688), .B(n1687), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[14])
         );
  OAI2BB1X1 U6759 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_3), 
        .B0(n2140), .Y(n2158) );
  AOI22X1 U6760 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_2), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[2]), 
        .B1(n17), .Y(n2140) );
  XOR2X1 U6761 ( .A(n1711), .B(n1712), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[2])
         );
  OAI2BB1X1 U6762 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_5), 
        .B0(n2138), .Y(n2156) );
  AOI22X1 U6763 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_4), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[4]), 
        .B1(n17), .Y(n2138) );
  XOR2X1 U6764 ( .A(n1707), .B(n1708), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[4])
         );
  OAI2BB1X1 U6765 ( .A0N(n368), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_7), 
        .B0(n2136), .Y(n2154) );
  AOI22X1 U6766 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_6), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[6]), 
        .B1(n17), .Y(n2136) );
  XOR2X1 U6767 ( .A(n1703), .B(n1704), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[6])
         );
  OAI2BB1X1 U6768 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_9), 
        .B0(n2134), .Y(n2152) );
  AOI22X1 U6769 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_8), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[8]), 
        .B1(n17), .Y(n2134) );
  XOR2X1 U6770 ( .A(n1699), .B(n1700), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[8])
         );
  OAI2BB1X1 U6771 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_11), 
        .B0(n2132), .Y(n2150) );
  AOI22X1 U6772 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_10), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[10]), 
        .B1(n17), .Y(n2132) );
  XOR2X1 U6773 ( .A(n1728), .B(n1727), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[10])
         );
  OAI2BB1X1 U6774 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_13), 
        .B0(n2130), .Y(n2148) );
  AOI22X1 U6775 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_12), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[12]), 
        .B1(n17), .Y(n2130) );
  XOR2X1 U6776 ( .A(n1724), .B(n1723), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[12])
         );
  OAI2BB1X1 U6777 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_15), 
        .B0(n2128), .Y(n2146) );
  AOI22X1 U6778 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_14), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[14]), 
        .B1(n17), .Y(n2128) );
  XOR2X1 U6779 ( .A(n1720), .B(n1719), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[14])
         );
  OAI2BB1X1 U6780 ( .A0N(n368), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_3), 
        .B0(n2249), .Y(n2267) );
  AOI22X1 U6781 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_2), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[2]), 
        .B1(n18), .Y(n2249) );
  XOR2X1 U6782 ( .A(n1743), .B(n1744), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[2])
         );
  OAI2BB1X1 U6783 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_5), 
        .B0(n2247), .Y(n2265) );
  AOI22X1 U6784 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_4), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[4]), 
        .B1(n18), .Y(n2247) );
  XOR2X1 U6785 ( .A(n1739), .B(n1740), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[4])
         );
  OAI2BB1X1 U6786 ( .A0N(n370), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_7), 
        .B0(n2245), .Y(n2263) );
  AOI22X1 U6787 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_6), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[6]), 
        .B1(n18), .Y(n2245) );
  XOR2X1 U6788 ( .A(n1735), .B(n1736), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[6])
         );
  OAI2BB1X1 U6789 ( .A0N(n370), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_9), 
        .B0(n2243), .Y(n2261) );
  AOI22X1 U6790 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_8), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[8]), 
        .B1(n18), .Y(n2243) );
  XOR2X1 U6791 ( .A(n1731), .B(n1732), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[8])
         );
  OAI2BB1X1 U6792 ( .A0N(n369), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_11), 
        .B0(n2241), .Y(n2259) );
  AOI22X1 U6793 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_10), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[10]), 
        .B1(n18), .Y(n2241) );
  XOR2X1 U6794 ( .A(n1760), .B(n1759), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[10])
         );
  OAI2BB1X1 U6795 ( .A0N(n368), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_13), 
        .B0(n2239), .Y(n2257) );
  AOI22X1 U6796 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_12), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[12]), 
        .B1(n18), .Y(n2239) );
  XOR2X1 U6797 ( .A(n1756), .B(n1755), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[12])
         );
  OAI2BB1X1 U6798 ( .A0N(n367), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_15), 
        .B0(n2237), .Y(n2255) );
  AOI22X1 U6799 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_14), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[14]), 
        .B1(n18), .Y(n2237) );
  XOR2X1 U6800 ( .A(n1752), .B(n1751), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[14])
         );
  OAI2BB1X1 U6801 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxcentral_parallel_output_0), 
        .B0(n1814), .Y(n1832) );
  AOI22X1 U6802 ( 
        .A0(input_times_b0_div_componentxUDxshifted_substraction_result_0), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxshifted_substraction_result_0), 
        .B1(n14), .Y(n1814) );
  OAI2BB1X1 U6803 ( .A0N(n368), 
        .A1N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_0), 
        .B0(n1924), .Y(n1942) );
  AOI22X1 U6804 ( 
        .A0(input_p1_times_b1_div_componentxUDxshifted_substraction_result_0), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxshifted_substraction_result_0), 
        .B1(n15), .Y(n1924) );
  OAI2BB1X1 U6805 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_0), 
        .B0(n2033), .Y(n2051) );
  AOI22X1 U6806 ( 
        .A0(input_p2_times_b2_div_componentxUDxshifted_substraction_result_0), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxshifted_substraction_result_0), 
        .B1(n16), .Y(n2033) );
  OAI2BB1X1 U6807 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_0), 
        .B0(n2143), .Y(n2161) );
  AOI22X1 U6808 ( 
        .A0(output_p1_times_a1_div_componentxUDxshifted_substraction_result_0), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxshifted_substraction_result_0), 
        .B1(n17), .Y(n2143) );
  OAI2BB1X1 U6809 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_0), 
        .B0(n2252), .Y(n2270) );
  AOI22X1 U6810 ( 
        .A0(output_p2_times_a2_div_componentxUDxshifted_substraction_result_0), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxshifted_substraction_result_0), 
        .B1(n18), .Y(n2252) );
  OAI2BB1X1 U6811 ( 
        .A0N(input_times_b0_div_componentxUDxcentral_parallel_output_17), 
        .A1N(n371), .B0(n1797), .Y(n1815) );
  AOI22X1 U6812 ( 
        .A0(input_times_b0_div_componentxUDxcentral_parallel_output_16), 
        .A1(n2), 
        .B0(input_times_b0_div_componentxUDxsubstraction_result_too_long[16]), 
        .B1(n14), .Y(n1797) );
  XOR2X1 U6813 ( .A(input_times_b0_div_componentxUDxactually_substractsxn24), 
        .B(input_times_b0_div_componentxUDxactually_substractsxn23), 
        .Y(input_times_b0_div_componentxUDxsubstraction_result_too_long[16])
         );
  XNOR2X1 U6814 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_16), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[16]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn24) );
  OAI2BB1X1 U6815 ( 
        .A0N(input_p1_times_b1_div_componentxUDxcentral_parallel_output_17), 
        .A1N(n367), .B0(n1907), .Y(n1925) );
  AOI22X1 U6816 ( 
        .A0(input_p1_times_b1_div_componentxUDxcentral_parallel_output_16), 
        .A1(n3), 
        .B0(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[16]), 
        .B1(n15), .Y(n1907) );
  XOR2X1 U6817 ( .A(n1652), .B(n1651), 
        .Y(input_p1_times_b1_div_componentxUDxsubstraction_result_too_long[16])
         );
  XNOR2X1 U6818 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_16), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[16]), 
        .Y(n1652) );
  OAI2BB1X1 U6819 ( 
        .A0N(input_p2_times_b2_div_componentxUDxcentral_parallel_output_17), 
        .A1N(n372), .B0(n2016), .Y(n2034) );
  AOI22X1 U6820 ( 
        .A0(input_p2_times_b2_div_componentxUDxcentral_parallel_output_16), 
        .A1(n4), 
        .B0(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[16]), 
        .B1(n16), .Y(n2016) );
  XOR2X1 U6821 ( .A(n1684), .B(n1683), 
        .Y(input_p2_times_b2_div_componentxUDxsubstraction_result_too_long[16])
         );
  XNOR2X1 U6822 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_16), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[16]), 
        .Y(n1684) );
  OAI2BB1X1 U6823 ( 
        .A0N(output_p1_times_a1_div_componentxUDxcentral_parallel_output_17), 
        .A1N(n370), .B0(n2126), .Y(n2144) );
  AOI22X1 U6824 ( 
        .A0(output_p1_times_a1_div_componentxUDxcentral_parallel_output_16), 
        .A1(n5), 
        .B0(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[16]), 
        .B1(n17), .Y(n2126) );
  XOR2X1 U6825 ( .A(n1716), .B(n1715), 
        .Y(output_p1_times_a1_div_componentxUDxsubstraction_result_too_long[16])
         );
  XNOR2X1 U6826 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_16), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[16]), 
        .Y(n1716) );
  OAI2BB1X1 U6827 ( 
        .A0N(output_p2_times_a2_div_componentxUDxcentral_parallel_output_17), 
        .A1N(n367), .B0(n2235), .Y(n2253) );
  AOI22X1 U6828 ( 
        .A0(output_p2_times_a2_div_componentxUDxcentral_parallel_output_16), 
        .A1(n6), 
        .B0(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[16]), 
        .B1(n18), .Y(n2235) );
  XOR2X1 U6829 ( .A(n1748), .B(n1747), 
        .Y(output_p2_times_a2_div_componentxUDxsubstraction_result_too_long[16])
         );
  XNOR2X1 U6830 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_16), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[16]), 
        .Y(n1748) );
  XOR2X1 U6831 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_5), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[5]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn10) );
  XOR2X1 U6832 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_5), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[5]), 
        .Y(n1642) );
  XOR2X1 U6833 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_5), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[5]), 
        .Y(n1674) );
  XOR2X1 U6834 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_5), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[5]), 
        .Y(n1706) );
  XOR2X1 U6835 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_5), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[5]), 
        .Y(n1738) );
  XOR2X1 U6836 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_7), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[7]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn6) );
  XOR2X1 U6837 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_7), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[7]), 
        .Y(n1638) );
  XOR2X1 U6838 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_7), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[7]), 
        .Y(n1670) );
  XOR2X1 U6839 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_7), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[7]), 
        .Y(n1702) );
  XOR2X1 U6840 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_7), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[7]), 
        .Y(n1734) );
  XNOR2X1 U6841 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_4), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[4]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn11) );
  XNOR2X1 U6842 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_4), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[4]), 
        .Y(n1643) );
  XNOR2X1 U6843 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_4), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[4]), 
        .Y(n1675) );
  XNOR2X1 U6844 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_4), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[4]), 
        .Y(n1707) );
  XNOR2X1 U6845 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_4), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[4]), 
        .Y(n1739) );
  XNOR2X1 U6846 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_6), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[6]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn7) );
  XNOR2X1 U6847 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_6), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[6]), 
        .Y(n1639) );
  XNOR2X1 U6848 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_6), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[6]), 
        .Y(n1671) );
  XNOR2X1 U6849 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_6), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[6]), 
        .Y(n1703) );
  XNOR2X1 U6850 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_6), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[6]), 
        .Y(n1735) );
  OAI2BB1X1 U6851 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[0]), 
        .B0(n1850), .Y(n1868) );
  NAND2X1 U6852 ( .A(n837), .B(en), .Y(n1850) );
  OAI2BB1X1 U6853 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[0]), 
        .B0(n1960), .Y(n1978) );
  NAND2X1 U6854 ( .A(n996), .B(en), .Y(n1960) );
  OAI2BB1X1 U6855 ( .A0N(n369), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[0]), 
        .B0(n2069), .Y(n2087) );
  NAND2X1 U6856 ( .A(n1155), .B(en), .Y(n2069) );
  OAI2BB1X1 U6857 ( .A0N(n369), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[0]), 
        .B0(n2179), .Y(n2197) );
  NAND2X1 U6858 ( .A(n519), .B(en), .Y(n2179) );
  OAI2BB1X1 U6859 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[0]), 
        .B0(n2288), .Y(n2306) );
  NAND2X1 U6860 ( .A(n678), .B(en), .Y(n2288) );
  XOR2X1 U6861 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_9), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[9]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn2) );
  XOR2X1 U6862 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_9), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[9]), 
        .Y(n1634) );
  XOR2X1 U6863 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_9), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[9]), 
        .Y(n1666) );
  XOR2X1 U6864 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_9), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[9]), 
        .Y(n1698) );
  XOR2X1 U6865 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_9), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[9]), 
        .Y(n1730) );
  XOR2X1 U6866 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_11), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[11]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn34) );
  XOR2X1 U6867 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_11), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[11]), 
        .Y(n1662) );
  XOR2X1 U6868 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_11), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[11]), 
        .Y(n1694) );
  XOR2X1 U6869 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_11), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[11]), 
        .Y(n1726) );
  XOR2X1 U6870 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_11), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[11]), 
        .Y(n1758) );
  XNOR2X1 U6871 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_8), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[8]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn3) );
  XNOR2X1 U6872 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_8), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[8]), 
        .Y(n1635) );
  XNOR2X1 U6873 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_8), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[8]), 
        .Y(n1667) );
  XNOR2X1 U6874 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_8), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[8]), 
        .Y(n1699) );
  XNOR2X1 U6875 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_8), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[8]), 
        .Y(n1731) );
  XNOR2X1 U6876 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_10), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[10]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn36) );
  XNOR2X1 U6877 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_10), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[10]), 
        .Y(n1664) );
  XNOR2X1 U6878 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_10), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[10]), 
        .Y(n1696) );
  XNOR2X1 U6879 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_10), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[10]), 
        .Y(n1728) );
  XNOR2X1 U6880 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_10), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[10]), 
        .Y(n1760) );
  XNOR2X1 U6881 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_12), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[12]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn32) );
  XNOR2X1 U6882 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_12), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[12]), 
        .Y(n1660) );
  XNOR2X1 U6883 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_12), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[12]), 
        .Y(n1692) );
  XNOR2X1 U6884 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_12), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[12]), 
        .Y(n1724) );
  XNOR2X1 U6885 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_12), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[12]), 
        .Y(n1756) );
  INVX1 U6886 ( .A(input_times_b0_div_componentxUDxcentral_parallel_output_9), 
        .Y(n1529) );
  INVX1 U6887 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_9), 
        .Y(n1513) );
  INVX1 U6888 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_9), 
        .Y(n1497) );
  INVX1 U6889 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_9), 
        .Y(n1481) );
  INVX1 U6890 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_9), 
        .Y(n1465) );
  BUFX4 U6891 ( .A(n4673), .Y(change_input) );
  XOR2X1 U6892 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_13), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[13]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn30) );
  XOR2X1 U6893 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_13), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[13]), 
        .Y(n1658) );
  XOR2X1 U6894 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_13), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[13]), 
        .Y(n1690) );
  XOR2X1 U6895 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_13), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[13]), 
        .Y(n1722) );
  XOR2X1 U6896 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_13), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[13]), 
        .Y(n1754) );
  XOR2X1 U6897 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_15), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[15]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn26) );
  XOR2X1 U6898 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_15), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[15]), 
        .Y(n1654) );
  XOR2X1 U6899 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_15), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[15]), 
        .Y(n1686) );
  XOR2X1 U6900 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_15), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[15]), 
        .Y(n1718) );
  XOR2X1 U6901 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_15), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[15]), 
        .Y(n1750) );
  XNOR2X1 U6902 ( 
        .A(input_times_b0_div_componentxUDxcentral_parallel_output_14), 
        .B(input_times_b0_div_componentxUDxsub_ready_negative_divisor[14]), 
        .Y(input_times_b0_div_componentxUDxactually_substractsxn28) );
  XNOR2X1 U6903 ( 
        .A(input_p1_times_b1_div_componentxUDxcentral_parallel_output_14), 
        .B(input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor[14]), 
        .Y(n1656) );
  XNOR2X1 U6904 ( 
        .A(input_p2_times_b2_div_componentxUDxcentral_parallel_output_14), 
        .B(input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor[14]), 
        .Y(n1688) );
  XNOR2X1 U6905 ( 
        .A(output_p1_times_a1_div_componentxUDxcentral_parallel_output_14), 
        .B(output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor[14]), 
        .Y(n1720) );
  XNOR2X1 U6906 ( 
        .A(output_p2_times_a2_div_componentxUDxcentral_parallel_output_14), 
        .B(output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor[14]), 
        .Y(n1752) );
  OAI2BB2X1 U6907 ( .B0(n1191), .B1(n321), .A0N(input_previous_1[9]), 
        .A1N(n321), .Y(n4628) );
  OAI2BB2X1 U6908 ( .B0(n1293), .B1(n1260), .A0N(input_previous_2[9]), 
        .A1N(n320), .Y(n4646) );
  OAI2BB2X1 U6909 ( .B0(n1198), .B1(n1260), .A0N(input_previous_1[16]), 
        .A1N(n321), .Y(n4635) );
  INVX1 U6910 ( .A(input_previous_0[16]), .Y(n1198) );
  OAI2BB2X1 U6911 ( .B0(n1197), .B1(n1260), .A0N(input_previous_1[15]), 
        .A1N(n321), .Y(n4634) );
  INVX1 U6912 ( .A(input_previous_0[15]), .Y(n1197) );
  OAI2BB2X1 U6913 ( .B0(n1196), .B1(n320), .A0N(input_previous_1[14]), 
        .A1N(n321), .Y(n4633) );
  INVX1 U6914 ( .A(input_previous_0[14]), .Y(n1196) );
  OAI2BB2X1 U6915 ( .B0(n1195), .B1(n1260), .A0N(input_previous_1[13]), 
        .A1N(n321), .Y(n4632) );
  INVX1 U6916 ( .A(input_previous_0[13]), .Y(n1195) );
  OAI2BB2X1 U6917 ( .B0(n1194), .B1(n1260), .A0N(input_previous_1[12]), 
        .A1N(n321), .Y(n4631) );
  INVX1 U6918 ( .A(input_previous_0[12]), .Y(n1194) );
  OAI2BB2X1 U6919 ( .B0(n1193), .B1(n319), .A0N(input_previous_1[11]), 
        .A1N(n321), .Y(n4630) );
  INVX1 U6920 ( .A(input_previous_0[11]), .Y(n1193) );
  OAI2BB2X1 U6921 ( .B0(n1192), .B1(n319), .A0N(input_previous_1[10]), 
        .A1N(n321), .Y(n4629) );
  INVX1 U6922 ( .A(input_previous_0[10]), .Y(n1192) );
  OAI2BB2X1 U6923 ( .B0(n1190), .B1(n1260), .A0N(input_previous_1[8]), 
        .A1N(n321), .Y(n4627) );
  INVX1 U6924 ( .A(input_previous_0[8]), .Y(n1190) );
  OAI2BB2X1 U6925 ( .B0(n1189), .B1(n1260), .A0N(input_previous_1[7]), 
        .A1N(n321), .Y(n4626) );
  INVX1 U6926 ( .A(input_previous_0[7]), .Y(n1189) );
  OAI2BB2X1 U6927 ( .B0(n1188), .B1(n1260), .A0N(input_previous_1[6]), 
        .A1N(n321), .Y(n4625) );
  INVX1 U6928 ( .A(input_previous_0[6]), .Y(n1188) );
  OAI2BB2X1 U6929 ( .B0(n1187), .B1(n321), .A0N(input_previous_1[5]), 
        .A1N(n321), .Y(n4624) );
  INVX1 U6930 ( .A(input_previous_0[5]), .Y(n1187) );
  OAI2BB2X1 U6931 ( .B0(n1186), .B1(n1260), .A0N(input_previous_1[4]), 
        .A1N(n321), .Y(n4623) );
  INVX1 U6932 ( .A(input_previous_0[4]), .Y(n1186) );
  OAI2BB2X1 U6933 ( .B0(n1185), .B1(n1260), .A0N(input_previous_1[3]), 
        .A1N(n321), .Y(n4622) );
  INVX1 U6934 ( .A(input_previous_0[3]), .Y(n1185) );
  OAI2BB2X1 U6935 ( .B0(n1184), .B1(n1260), .A0N(input_previous_1[2]), 
        .A1N(n321), .Y(n4621) );
  INVX1 U6936 ( .A(input_previous_0[2]), .Y(n1184) );
  OAI2BB2X1 U6937 ( .B0(n1183), .B1(n321), .A0N(input_previous_1[1]), 
        .A1N(n321), .Y(n4620) );
  INVX1 U6938 ( .A(input_previous_0[1]), .Y(n1183) );
  OAI2BB2X1 U6939 ( .B0(n1182), .B1(n1260), 
        .A0N(input_p1_times_b1_mul_componentxinput_A_inverted[0]), .A1N(n319), 
        .Y(n4619) );
  INVX1 U6940 ( .A(input_times_b0_mul_componentxinput_A_inverted[0]), 
        .Y(n1182) );
  OAI2BB2X1 U6941 ( .B0(n1300), .B1(n1260), .A0N(input_previous_2[16]), 
        .A1N(n320), .Y(n4653) );
  INVX1 U6942 ( .A(input_previous_1[16]), .Y(n1300) );
  OAI2BB2X1 U6943 ( .B0(n1299), .B1(n1260), .A0N(input_previous_2[15]), 
        .A1N(n320), .Y(n4652) );
  INVX1 U6944 ( .A(input_previous_1[15]), .Y(n1299) );
  OAI2BB2X1 U6945 ( .B0(n1298), .B1(n1260), .A0N(input_previous_2[14]), 
        .A1N(n320), .Y(n4651) );
  INVX1 U6946 ( .A(input_previous_1[14]), .Y(n1298) );
  OAI2BB2X1 U6947 ( .B0(n1297), .B1(n321), .A0N(input_previous_2[13]), 
        .A1N(n320), .Y(n4650) );
  INVX1 U6948 ( .A(input_previous_1[13]), .Y(n1297) );
  OAI2BB2X1 U6949 ( .B0(n1296), .B1(n1260), .A0N(input_previous_2[12]), 
        .A1N(n320), .Y(n4649) );
  INVX1 U6950 ( .A(input_previous_1[12]), .Y(n1296) );
  OAI2BB2X1 U6951 ( .B0(n1295), .B1(n1260), .A0N(input_previous_2[11]), 
        .A1N(n320), .Y(n4648) );
  INVX1 U6952 ( .A(input_previous_1[11]), .Y(n1295) );
  OAI2BB2X1 U6953 ( .B0(n1294), .B1(n320), .A0N(input_previous_2[10]), 
        .A1N(n320), .Y(n4647) );
  INVX1 U6954 ( .A(input_previous_1[10]), .Y(n1294) );
  OAI2BB2X1 U6955 ( .B0(n1292), .B1(n1260), .A0N(input_previous_2[8]), 
        .A1N(n320), .Y(n4645) );
  INVX1 U6956 ( .A(input_previous_1[8]), .Y(n1292) );
  OAI2BB2X1 U6957 ( .B0(n1291), .B1(n319), .A0N(input_previous_2[7]), 
        .A1N(n320), .Y(n4644) );
  INVX1 U6958 ( .A(input_previous_1[7]), .Y(n1291) );
  OAI2BB2X1 U6959 ( .B0(n1290), .B1(n321), .A0N(input_previous_2[6]), 
        .A1N(n321), .Y(n4643) );
  INVX1 U6960 ( .A(input_previous_1[6]), .Y(n1290) );
  OAI2BB2X1 U6961 ( .B0(n1289), .B1(n320), .A0N(input_previous_2[5]), 
        .A1N(n321), .Y(n4642) );
  INVX1 U6962 ( .A(input_previous_1[5]), .Y(n1289) );
  OAI2BB2X1 U6963 ( .B0(n1288), .B1(n319), .A0N(input_previous_2[4]), 
        .A1N(n321), .Y(n4641) );
  INVX1 U6964 ( .A(input_previous_1[4]), .Y(n1288) );
  OAI2BB2X1 U6965 ( .B0(n1287), .B1(n321), .A0N(input_previous_2[3]), 
        .A1N(n321), .Y(n4640) );
  INVX1 U6966 ( .A(input_previous_1[3]), .Y(n1287) );
  OAI2BB2X1 U6967 ( .B0(n1286), .B1(n320), .A0N(input_previous_2[2]), 
        .A1N(n321), .Y(n4639) );
  INVX1 U6968 ( .A(input_previous_1[2]), .Y(n1286) );
  OAI2BB2X1 U6969 ( .B0(n1285), .B1(n320), .A0N(input_previous_2[1]), 
        .A1N(n321), .Y(n4638) );
  INVX1 U6970 ( .A(input_previous_1[1]), .Y(n1285) );
  OAI2BB2X1 U6971 ( .B0(n1284), .B1(n319), 
        .A0N(input_p2_times_b2_mul_componentxinput_A_inverted[0]), .A1N(n321), 
        .Y(n4637) );
  INVX1 U6972 ( .A(input_p1_times_b1_mul_componentxinput_A_inverted[0]), 
        .Y(n1284) );
  OAI2BB2X1 U6973 ( .B0(n1174), .B1(n320), .A0N(input_previous_0[16]), 
        .A1N(n319), .Y(input_prev_0_registerxn18) );
  OAI2BB2X1 U6974 ( .B0(n1174), .B1(n321), .A0N(input_previous_0[15]), 
        .A1N(n320), .Y(input_prev_0_registerxn17) );
  OAI2BB2X1 U6975 ( .B0(n1174), .B1(n1260), .A0N(input_previous_0[14]), 
        .A1N(n319), .Y(input_prev_0_registerxn16) );
  OAI2BB2X1 U6976 ( .B0(n1174), .B1(n321), .A0N(input_previous_0[13]), 
        .A1N(n319), .Y(input_prev_0_registerxn15) );
  OAI2BB2X1 U6977 ( .B0(n1174), .B1(n1260), .A0N(input_previous_0[12]), 
        .A1N(n319), .Y(input_prev_0_registerxn14) );
  OAI2BB2X1 U6978 ( .B0(n1174), .B1(n1260), .A0N(input_previous_0[11]), 
        .A1N(n319), .Y(input_prev_0_registerxn13) );
  OAI2BB2X1 U6979 ( .B0(n1174), .B1(n320), .A0N(input_previous_0[10]), 
        .A1N(n319), .Y(input_prev_0_registerxn12) );
  OAI2BB2X1 U6980 ( .B0(n1174), .B1(n1260), .A0N(input_previous_0[9]), 
        .A1N(n319), .Y(input_prev_0_registerxn11) );
  OAI2BB2X1 U6981 ( .B0(n1174), .B1(n321), .A0N(input_previous_0[8]), 
        .A1N(n319), .Y(input_prev_0_registerxn10) );
  OAI2BB2X1 U6982 ( .B0(n1174), .B1(n320), .A0N(input_previous_0[7]), 
        .A1N(n319), .Y(input_prev_0_registerxn9) );
  OAI2BB2X1 U6983 ( .B0(n1175), .B1(n319), .A0N(input_previous_0[6]), 
        .A1N(n319), .Y(input_prev_0_registerxn8) );
  INVX1 U6984 ( .A(\input_signal[6] ), .Y(n1175) );
  OAI2BB2X1 U6985 ( .B0(n1176), .B1(n1260), .A0N(input_previous_0[5]), 
        .A1N(n319), .Y(input_prev_0_registerxn7) );
  INVX1 U6986 ( .A(\input_signal[5] ), .Y(n1176) );
  OAI2BB2X1 U6987 ( .B0(n1177), .B1(n1260), .A0N(input_previous_0[4]), 
        .A1N(n319), .Y(input_prev_0_registerxn6) );
  INVX1 U6988 ( .A(\input_signal[4] ), .Y(n1177) );
  OAI2BB2X1 U6989 ( .B0(n1178), .B1(n321), .A0N(input_previous_0[3]), 
        .A1N(n319), .Y(input_prev_0_registerxn5) );
  INVX1 U6990 ( .A(\input_signal[3] ), .Y(n1178) );
  OAI2BB2X1 U6991 ( .B0(n1179), .B1(n1260), .A0N(input_previous_0[2]), 
        .A1N(n319), .Y(input_prev_0_registerxn4) );
  INVX1 U6992 ( .A(\input_signal[2] ), .Y(n1179) );
  OAI2BB2X1 U6993 ( .B0(n1180), .B1(n319), .A0N(input_previous_0[1]), 
        .A1N(n319), .Y(input_prev_0_registerxn3) );
  INVX1 U6994 ( .A(\input_signal[1] ), .Y(n1180) );
  OAI2BB2X1 U6995 ( .B0(n1181), .B1(n1260), 
        .A0N(input_times_b0_mul_componentxinput_A_inverted[0]), .A1N(n319), 
        .Y(input_prev_0_registerxn2) );
  INVX1 U6996 ( .A(\input_signal[0] ), .Y(n1181) );
  NAND2X1 U6997 ( .A(change_input), .B(en), .Y(n109) );
  INVX1 U6998 ( .A(n109), .Y(n1871) );
  NAND2X1 U6999 ( .A(change_input), .B(en), .Y(n110) );
  INVX1 U7000 ( .A(n110), .Y(n2090) );
  NAND2X1 U7001 ( .A(input_p1_times_b1_div_componentxoutput_ready_signal), 
        .B(en), .Y(n4203) );
  NAND2X1 U7002 ( .A(input_p2_times_b2_div_componentxoutput_ready_signal), 
        .B(en), .Y(n4259) );
  NAND2X1 U7003 ( .A(n7), .B(en), .Y(n4369) );
  NAND2X1 U7004 ( .A(n8), .B(en), .Y(input_times_b0_div_componentxn24) );
  OAI22X1 U7005 ( .A0(n374), .A1(n151), .B0(n1381), .B1(n4203), .Y(n4240) );
  INVX1 U7006 ( .A(input_p1_times_b1_div_componentxoutput_sign_gated_prev), 
        .Y(n1381) );
  OAI22X1 U7007 ( .A0(n376), .A1(n149), .B0(n1361), .B1(n4259), .Y(n4296) );
  INVX1 U7008 ( .A(input_p2_times_b2_div_componentxoutput_sign_gated_prev), 
        .Y(n1361) );
  OAI22X1 U7009 ( .A0(n378), .A1(n145), .B0(n1322), .B1(n4369), .Y(n4406) );
  INVX1 U7010 ( .A(output_p2_times_a2_div_componentxoutput_sign_gated_prev), 
        .Y(n1322) );
  OAI22X1 U7011 ( .A0(n380), .A1(n135), .B0(n1239), 
        .B1(input_times_b0_div_componentxn24), 
        .Y(input_times_b0_div_componentxn62) );
  INVX1 U7012 ( .A(input_times_b0_div_componentxoutput_sign_gated_prev), 
        .Y(n1239) );
  OAI22X1 U7013 ( .A0(n367), .A1(n1252), .B0(en), .B1(n1251), 
        .Y(clock_chopper_and_divisionxn37) );
  OAI22X1 U7014 ( .A0(en), .A1(n1240), .B0(n1241), .B1(n367), 
        .Y(clock_chopper_and_divisionxn26) );
  OAI22X1 U7015 ( .A0(en), .A1(n1259), .B0(n367), .B1(n1261), 
        .Y(clock_chopper_and_divisionxn45) );
  OAI22X1 U7016 ( .A0(en), .A1(n1258), .B0(n368), .B1(n1259), 
        .Y(clock_chopper_and_divisionxn44) );
  OAI22X1 U7017 ( .A0(en), .A1(n1257), .B0(n367), .B1(n1258), 
        .Y(clock_chopper_and_divisionxn43) );
  OAI22X1 U7018 ( .A0(en), .A1(n1256), .B0(n367), .B1(n1257), 
        .Y(clock_chopper_and_divisionxn42) );
  OAI22X1 U7019 ( .A0(en), .A1(n1255), .B0(n367), .B1(n1256), 
        .Y(clock_chopper_and_divisionxn41) );
  OAI22X1 U7020 ( .A0(en), .A1(n1254), .B0(n370), .B1(n1255), 
        .Y(clock_chopper_and_divisionxn40) );
  OAI22X1 U7021 ( .A0(en), .A1(n1253), .B0(n367), .B1(n1254), 
        .Y(clock_chopper_and_divisionxn39) );
  OAI22X1 U7022 ( .A0(en), .A1(n1252), .B0(n369), .B1(n1253), 
        .Y(clock_chopper_and_divisionxn38) );
  OAI22X1 U7023 ( .A0(en), .A1(n1250), .B0(n368), .B1(n1251), 
        .Y(clock_chopper_and_divisionxn36) );
  OAI22X1 U7024 ( .A0(en), .A1(n1249), .B0(n367), .B1(n1250), 
        .Y(clock_chopper_and_divisionxn35) );
  OAI22X1 U7025 ( .A0(en), .A1(n1248), .B0(n369), .B1(n1249), 
        .Y(clock_chopper_and_divisionxn34) );
  OAI22X1 U7026 ( .A0(en), .A1(n1247), .B0(n368), .B1(n1248), 
        .Y(clock_chopper_and_divisionxn33) );
  OAI22X1 U7027 ( .A0(en), .A1(n1246), .B0(n367), .B1(n1247), 
        .Y(clock_chopper_and_divisionxn32) );
  OAI22X1 U7028 ( .A0(en), .A1(n1245), .B0(n367), .B1(n1246), 
        .Y(clock_chopper_and_divisionxn31) );
  OAI22X1 U7029 ( .A0(en), .A1(n1244), .B0(n367), .B1(n1245), 
        .Y(clock_chopper_and_divisionxn30) );
  OAI22X1 U7030 ( .A0(en), .A1(n1243), .B0(n367), .B1(n1244), 
        .Y(clock_chopper_and_divisionxn29) );
  OAI22X1 U7031 ( .A0(en), .A1(n1242), .B0(n367), .B1(n1243), 
        .Y(clock_chopper_and_divisionxn28) );
  OAI22X1 U7032 ( .A0(en), .A1(n1241), .B0(n367), .B1(n1242), 
        .Y(clock_chopper_and_divisionxn27) );
  OAI22X1 U7033 ( .A0(n367), .A1(n1240), .B0(en), .B1(n1262), 
        .Y(clock_chopper_and_divisionxn49) );
  OAI22X1 U7034 ( .A0(en), .A1(n1261), .B0(n367), .B1(n1262), 
        .Y(clock_chopper_and_divisionxn47) );
  INVX1 U7035 ( .A(input_p1_times_b1_div_componentxoutput_ready_signal), 
        .Y(n161) );
  INVX1 U7036 ( .A(input_p2_times_b2_div_componentxoutput_ready_signal), 
        .Y(n162) );
  INVX1 U7037 ( .A(output_p1_times_a1_div_componentxoutput_ready_signal), 
        .Y(n163) );
  OAI2BB2X1 U7038 ( .B0(n367), .B1(n1261), .A0N(n258), .A1N(n368), 
        .Y(clock_chopper_and_divisionxn46) );
  BUFX3 U7039 ( .A(n4673), .Y(n258) );
  INVX1 U7040 ( .A(clock_chopper_and_divisionxdivision_ring[20]), .Y(n1241) );
  INVX1 U7041 ( .A(clock_chopper_and_divisionxdivision_ring[9]), .Y(n1252) );
  INVX1 U7042 ( .A(clock_chopper_and_divisionxdivision_ring[21]), .Y(n1240) );
  INVX1 U7043 ( .A(clock_chopper_and_divisionxdivision_ring[2]), .Y(n1259) );
  INVX1 U7044 ( .A(clock_chopper_and_divisionxdivision_ring[3]), .Y(n1258) );
  INVX1 U7045 ( .A(clock_chopper_and_divisionxdivision_ring[4]), .Y(n1257) );
  INVX1 U7046 ( .A(clock_chopper_and_divisionxdivision_ring[5]), .Y(n1256) );
  INVX1 U7047 ( .A(clock_chopper_and_divisionxdivision_ring[6]), .Y(n1255) );
  INVX1 U7048 ( .A(clock_chopper_and_divisionxdivision_ring[7]), .Y(n1254) );
  INVX1 U7049 ( .A(clock_chopper_and_divisionxdivision_ring[8]), .Y(n1253) );
  INVX1 U7050 ( .A(clock_chopper_and_divisionxdivision_ring[11]), .Y(n1250) );
  INVX1 U7051 ( .A(clock_chopper_and_divisionxdivision_ring[12]), .Y(n1249) );
  INVX1 U7052 ( .A(clock_chopper_and_divisionxdivision_ring[13]), .Y(n1248) );
  INVX1 U7053 ( .A(clock_chopper_and_divisionxdivision_ring[14]), .Y(n1247) );
  INVX1 U7054 ( .A(clock_chopper_and_divisionxdivision_ring[15]), .Y(n1246) );
  INVX1 U7055 ( .A(clock_chopper_and_divisionxdivision_ring[16]), .Y(n1245) );
  INVX1 U7056 ( .A(clock_chopper_and_divisionxdivision_ring[17]), .Y(n1244) );
  INVX1 U7057 ( .A(clock_chopper_and_divisionxdivision_ring[18]), .Y(n1243) );
  INVX1 U7058 ( .A(clock_chopper_and_divisionxdivision_ring[19]), .Y(n1242) );
  INVX1 U7059 ( .A(clock_chopper_and_divisionxdivision_ring[10]), .Y(n1251) );
  OAI2BB1X1 U7060 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[1]), 
        .B0(n1849), .Y(n1867) );
  NAND2X1 U7061 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[0]), 
        .B(en), .Y(n1849) );
  OAI2BB1X1 U7062 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[2]), 
        .B0(n1848), .Y(n1866) );
  NAND2X1 U7063 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[1]), 
        .B(en), .Y(n1848) );
  OAI2BB1X1 U7064 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[3]), 
        .B0(n1847), .Y(n1865) );
  NAND2X1 U7065 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[2]), 
        .B(en), .Y(n1847) );
  OAI2BB1X1 U7066 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[4]), 
        .B0(n1846), .Y(n1864) );
  NAND2X1 U7067 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[3]), 
        .B(en), .Y(n1846) );
  OAI2BB1X1 U7068 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[5]), 
        .B0(n1845), .Y(n1863) );
  NAND2X1 U7069 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[4]), 
        .B(en), .Y(n1845) );
  OAI2BB1X1 U7070 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[6]), 
        .B0(n1844), .Y(n1862) );
  NAND2X1 U7071 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[5]), 
        .B(en), .Y(n1844) );
  OAI2BB1X1 U7072 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[7]), 
        .B0(n1843), .Y(n1861) );
  NAND2X1 U7073 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[6]), 
        .B(en), .Y(n1843) );
  OAI2BB1X1 U7074 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[8]), 
        .B0(n1842), .Y(n1860) );
  NAND2X1 U7075 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[7]), 
        .B(en), .Y(n1842) );
  OAI2BB1X1 U7076 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[9]), 
        .B0(n1841), .Y(n1859) );
  NAND2X1 U7077 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[8]), 
        .B(en), .Y(n1841) );
  OAI2BB1X1 U7078 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[10]), 
        .B0(n1840), .Y(n1858) );
  NAND2X1 U7079 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[9]), 
        .B(en), .Y(n1840) );
  OAI2BB1X1 U7080 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[11]), 
        .B0(n1839), .Y(n1857) );
  NAND2X1 U7081 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[10]), 
        .B(en), .Y(n1839) );
  OAI2BB1X1 U7082 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[12]), 
        .B0(n1838), .Y(n1856) );
  NAND2X1 U7083 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[11]), 
        .B(en), .Y(n1838) );
  OAI2BB1X1 U7084 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[13]), 
        .B0(n1837), .Y(n1855) );
  NAND2X1 U7085 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[12]), 
        .B(en), .Y(n1837) );
  OAI2BB1X1 U7086 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[14]), 
        .B0(n1836), .Y(n1854) );
  NAND2X1 U7087 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[13]), 
        .B(en), .Y(n1836) );
  OAI2BB1X1 U7088 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[15]), 
        .B0(n1835), .Y(n1853) );
  NAND2X1 U7089 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[14]), 
        .B(en), .Y(n1835) );
  OAI2BB1X1 U7090 ( .A0N(n370), 
        .A1N(input_times_b0_div_componentxUDxquotient_not_gated[16]), 
        .B0(n1834), .Y(n1852) );
  NAND2X1 U7091 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[15]), 
        .B(en), .Y(n1834) );
  OAI2BB1X1 U7092 ( 
        .A0N(input_times_b0_div_componentxUDxquotient_not_gated[17]), 
        .A1N(n370), .B0(n1833), .Y(n1851) );
  NAND2X1 U7093 ( .A(input_times_b0_div_componentxUDxquotient_not_gated[16]), 
        .B(en), .Y(n1833) );
  OAI2BB1X1 U7094 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[1]), 
        .B0(n1959), .Y(n1977) );
  NAND2X1 U7095 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[0]), 
        .B(en), .Y(n1959) );
  OAI2BB1X1 U7096 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[2]), 
        .B0(n1958), .Y(n1976) );
  NAND2X1 U7097 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[1]), 
        .B(en), .Y(n1958) );
  OAI2BB1X1 U7098 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[3]), 
        .B0(n1957), .Y(n1975) );
  NAND2X1 U7099 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[2]), 
        .B(en), .Y(n1957) );
  OAI2BB1X1 U7100 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[4]), 
        .B0(n1956), .Y(n1974) );
  NAND2X1 U7101 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[3]), 
        .B(en), .Y(n1956) );
  OAI2BB1X1 U7102 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[5]), 
        .B0(n1955), .Y(n1973) );
  NAND2X1 U7103 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[4]), 
        .B(en), .Y(n1955) );
  OAI2BB1X1 U7104 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[6]), 
        .B0(n1954), .Y(n1972) );
  NAND2X1 U7105 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[5]), 
        .B(en), .Y(n1954) );
  OAI2BB1X1 U7106 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[7]), 
        .B0(n1953), .Y(n1971) );
  NAND2X1 U7107 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[6]), 
        .B(en), .Y(n1953) );
  OAI2BB1X1 U7108 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[8]), 
        .B0(n1952), .Y(n1970) );
  NAND2X1 U7109 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[7]), 
        .B(en), .Y(n1952) );
  OAI2BB1X1 U7110 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[9]), 
        .B0(n1951), .Y(n1969) );
  NAND2X1 U7111 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[8]), 
        .B(en), .Y(n1951) );
  OAI2BB1X1 U7112 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[10]), 
        .B0(n1950), .Y(n1968) );
  NAND2X1 U7113 ( .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[9]), 
        .B(en), .Y(n1950) );
  OAI2BB1X1 U7114 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[11]), 
        .B0(n1949), .Y(n1967) );
  NAND2X1 U7115 ( 
        .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[10]), .B(en), 
        .Y(n1949) );
  OAI2BB1X1 U7116 ( .A0N(n372), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[12]), 
        .B0(n1948), .Y(n1966) );
  NAND2X1 U7117 ( 
        .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[11]), .B(en), 
        .Y(n1948) );
  OAI2BB1X1 U7118 ( .A0N(n369), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[13]), 
        .B0(n1947), .Y(n1965) );
  NAND2X1 U7119 ( 
        .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[12]), .B(en), 
        .Y(n1947) );
  OAI2BB1X1 U7120 ( .A0N(n370), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[14]), 
        .B0(n1946), .Y(n1964) );
  NAND2X1 U7121 ( 
        .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[13]), .B(en), 
        .Y(n1946) );
  OAI2BB1X1 U7122 ( .A0N(n367), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[15]), 
        .B0(n1945), .Y(n1963) );
  NAND2X1 U7123 ( 
        .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[14]), .B(en), 
        .Y(n1945) );
  OAI2BB1X1 U7124 ( .A0N(n371), 
        .A1N(input_p1_times_b1_div_componentxUDxquotient_not_gated[16]), 
        .B0(n1944), .Y(n1962) );
  NAND2X1 U7125 ( 
        .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[15]), .B(en), 
        .Y(n1944) );
  OAI2BB1X1 U7126 ( 
        .A0N(input_p1_times_b1_div_componentxUDxquotient_not_gated[17]), 
        .A1N(n369), .B0(n1943), .Y(n1961) );
  NAND2X1 U7127 ( 
        .A(input_p1_times_b1_div_componentxUDxquotient_not_gated[16]), .B(en), 
        .Y(n1943) );
  OAI2BB1X1 U7128 ( .A0N(n372), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[1]), 
        .B0(n2068), .Y(n2086) );
  NAND2X1 U7129 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[0]), 
        .B(en), .Y(n2068) );
  OAI2BB1X1 U7130 ( .A0N(n371), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[2]), 
        .B0(n2067), .Y(n2085) );
  NAND2X1 U7131 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[1]), 
        .B(en), .Y(n2067) );
  OAI2BB1X1 U7132 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[3]), 
        .B0(n2066), .Y(n2084) );
  NAND2X1 U7133 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[2]), 
        .B(en), .Y(n2066) );
  OAI2BB1X1 U7134 ( .A0N(n367), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[4]), 
        .B0(n2065), .Y(n2083) );
  NAND2X1 U7135 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[3]), 
        .B(en), .Y(n2065) );
  OAI2BB1X1 U7136 ( .A0N(n372), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[5]), 
        .B0(n2064), .Y(n2082) );
  NAND2X1 U7137 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[4]), 
        .B(en), .Y(n2064) );
  OAI2BB1X1 U7138 ( .A0N(n371), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[6]), 
        .B0(n2063), .Y(n2081) );
  NAND2X1 U7139 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[5]), 
        .B(en), .Y(n2063) );
  OAI2BB1X1 U7140 ( .A0N(n371), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[7]), 
        .B0(n2062), .Y(n2080) );
  NAND2X1 U7141 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[6]), 
        .B(en), .Y(n2062) );
  OAI2BB1X1 U7142 ( .A0N(n371), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[8]), 
        .B0(n2061), .Y(n2079) );
  NAND2X1 U7143 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[7]), 
        .B(en), .Y(n2061) );
  OAI2BB1X1 U7144 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[9]), 
        .B0(n2060), .Y(n2078) );
  NAND2X1 U7145 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[8]), 
        .B(en), .Y(n2060) );
  OAI2BB1X1 U7146 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[10]), 
        .B0(n2059), .Y(n2077) );
  NAND2X1 U7147 ( .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[9]), 
        .B(en), .Y(n2059) );
  OAI2BB1X1 U7148 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[11]), 
        .B0(n2058), .Y(n2076) );
  NAND2X1 U7149 ( 
        .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[10]), .B(en), 
        .Y(n2058) );
  OAI2BB1X1 U7150 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[12]), 
        .B0(n2057), .Y(n2075) );
  NAND2X1 U7151 ( 
        .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[11]), .B(en), 
        .Y(n2057) );
  OAI2BB1X1 U7152 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[13]), 
        .B0(n2056), .Y(n2074) );
  NAND2X1 U7153 ( 
        .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[12]), .B(en), 
        .Y(n2056) );
  OAI2BB1X1 U7154 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[14]), 
        .B0(n2055), .Y(n2073) );
  NAND2X1 U7155 ( 
        .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[13]), .B(en), 
        .Y(n2055) );
  OAI2BB1X1 U7156 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[15]), 
        .B0(n2054), .Y(n2072) );
  NAND2X1 U7157 ( 
        .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[14]), .B(en), 
        .Y(n2054) );
  OAI2BB1X1 U7158 ( .A0N(n368), 
        .A1N(input_p2_times_b2_div_componentxUDxquotient_not_gated[16]), 
        .B0(n2053), .Y(n2071) );
  NAND2X1 U7159 ( 
        .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[15]), .B(en), 
        .Y(n2053) );
  OAI2BB1X1 U7160 ( 
        .A0N(input_p2_times_b2_div_componentxUDxquotient_not_gated[17]), 
        .A1N(n369), .B0(n2052), .Y(n2070) );
  NAND2X1 U7161 ( 
        .A(input_p2_times_b2_div_componentxUDxquotient_not_gated[16]), .B(en), 
        .Y(n2052) );
  OAI2BB1X1 U7162 ( .A0N(n371), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[1]), 
        .B0(n2178), .Y(n2196) );
  NAND2X1 U7163 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[0]), .B(en), 
        .Y(n2178) );
  OAI2BB1X1 U7164 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[2]), 
        .B0(n2177), .Y(n2195) );
  NAND2X1 U7165 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[1]), .B(en), 
        .Y(n2177) );
  OAI2BB1X1 U7166 ( .A0N(n370), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[3]), 
        .B0(n2176), .Y(n2194) );
  NAND2X1 U7167 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[2]), .B(en), 
        .Y(n2176) );
  OAI2BB1X1 U7168 ( .A0N(n367), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[4]), 
        .B0(n2175), .Y(n2193) );
  NAND2X1 U7169 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[3]), .B(en), 
        .Y(n2175) );
  OAI2BB1X1 U7170 ( .A0N(n368), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[5]), 
        .B0(n2174), .Y(n2192) );
  NAND2X1 U7171 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[4]), .B(en), 
        .Y(n2174) );
  OAI2BB1X1 U7172 ( .A0N(n369), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[6]), 
        .B0(n2173), .Y(n2191) );
  NAND2X1 U7173 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[5]), .B(en), 
        .Y(n2173) );
  OAI2BB1X1 U7174 ( .A0N(n371), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[7]), 
        .B0(n2172), .Y(n2190) );
  NAND2X1 U7175 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[6]), .B(en), 
        .Y(n2172) );
  OAI2BB1X1 U7176 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[8]), 
        .B0(n2171), .Y(n2189) );
  NAND2X1 U7177 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[7]), .B(en), 
        .Y(n2171) );
  OAI2BB1X1 U7178 ( .A0N(n370), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[9]), 
        .B0(n2170), .Y(n2188) );
  NAND2X1 U7179 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[8]), .B(en), 
        .Y(n2170) );
  OAI2BB1X1 U7180 ( .A0N(n367), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[10]), 
        .B0(n2169), .Y(n2187) );
  NAND2X1 U7181 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[9]), .B(en), 
        .Y(n2169) );
  OAI2BB1X1 U7182 ( .A0N(n368), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[11]), 
        .B0(n2168), .Y(n2186) );
  NAND2X1 U7183 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[10]), .B(en), 
        .Y(n2168) );
  OAI2BB1X1 U7184 ( .A0N(n369), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[12]), 
        .B0(n2167), .Y(n2185) );
  NAND2X1 U7185 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[11]), .B(en), 
        .Y(n2167) );
  OAI2BB1X1 U7186 ( .A0N(n371), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[13]), 
        .B0(n2166), .Y(n2184) );
  NAND2X1 U7187 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[12]), .B(en), 
        .Y(n2166) );
  OAI2BB1X1 U7188 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[14]), 
        .B0(n2165), .Y(n2183) );
  NAND2X1 U7189 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[13]), .B(en), 
        .Y(n2165) );
  OAI2BB1X1 U7190 ( .A0N(n372), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[15]), 
        .B0(n2164), .Y(n2182) );
  NAND2X1 U7191 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[14]), .B(en), 
        .Y(n2164) );
  OAI2BB1X1 U7192 ( .A0N(n370), 
        .A1N(output_p1_times_a1_div_componentxUDxquotient_not_gated[16]), 
        .B0(n2163), .Y(n2181) );
  NAND2X1 U7193 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[15]), .B(en), 
        .Y(n2163) );
  OAI2BB1X1 U7194 ( 
        .A0N(output_p1_times_a1_div_componentxUDxquotient_not_gated[17]), 
        .A1N(n368), .B0(n2162), .Y(n2180) );
  NAND2X1 U7195 ( 
        .A(output_p1_times_a1_div_componentxUDxquotient_not_gated[16]), .B(en), 
        .Y(n2162) );
  OAI2BB1X1 U7196 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[1]), 
        .B0(n2287), .Y(n2305) );
  NAND2X1 U7197 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[0]), .B(en), 
        .Y(n2287) );
  OAI2BB1X1 U7198 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[2]), 
        .B0(n2286), .Y(n2304) );
  NAND2X1 U7199 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[1]), .B(en), 
        .Y(n2286) );
  OAI2BB1X1 U7200 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[3]), 
        .B0(n2285), .Y(n2303) );
  NAND2X1 U7201 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[2]), .B(en), 
        .Y(n2285) );
  OAI2BB1X1 U7202 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[4]), 
        .B0(n2284), .Y(n2302) );
  NAND2X1 U7203 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[3]), .B(en), 
        .Y(n2284) );
  OAI2BB1X1 U7204 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[5]), 
        .B0(n2283), .Y(n2301) );
  NAND2X1 U7205 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[4]), .B(en), 
        .Y(n2283) );
  OAI2BB1X1 U7206 ( .A0N(n368), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[6]), 
        .B0(n2282), .Y(n2300) );
  NAND2X1 U7207 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[5]), .B(en), 
        .Y(n2282) );
  OAI2BB1X1 U7208 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[7]), 
        .B0(n2281), .Y(n2299) );
  NAND2X1 U7209 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[6]), .B(en), 
        .Y(n2281) );
  OAI2BB1X1 U7210 ( .A0N(n367), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[8]), 
        .B0(n2280), .Y(n2298) );
  NAND2X1 U7211 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[7]), .B(en), 
        .Y(n2280) );
  OAI2BB1X1 U7212 ( .A0N(n370), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[9]), 
        .B0(n2279), .Y(n2297) );
  NAND2X1 U7213 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[8]), .B(en), 
        .Y(n2279) );
  OAI2BB1X1 U7214 ( .A0N(n369), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[10]), 
        .B0(n2278), .Y(n2296) );
  NAND2X1 U7215 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[9]), .B(en), 
        .Y(n2278) );
  OAI2BB1X1 U7216 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[11]), 
        .B0(n2277), .Y(n2295) );
  NAND2X1 U7217 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[10]), .B(en), 
        .Y(n2277) );
  OAI2BB1X1 U7218 ( .A0N(n367), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[12]), 
        .B0(n2276), .Y(n2294) );
  NAND2X1 U7219 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[11]), .B(en), 
        .Y(n2276) );
  OAI2BB1X1 U7220 ( .A0N(n371), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[13]), 
        .B0(n2275), .Y(n2293) );
  NAND2X1 U7221 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[12]), .B(en), 
        .Y(n2275) );
  OAI2BB1X1 U7222 ( .A0N(n368), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[14]), 
        .B0(n2274), .Y(n2292) );
  NAND2X1 U7223 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[13]), .B(en), 
        .Y(n2274) );
  OAI2BB1X1 U7224 ( .A0N(n372), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[15]), 
        .B0(n2273), .Y(n2291) );
  NAND2X1 U7225 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[14]), .B(en), 
        .Y(n2273) );
  OAI2BB1X1 U7226 ( .A0N(n368), 
        .A1N(output_p2_times_a2_div_componentxUDxquotient_not_gated[16]), 
        .B0(n2272), .Y(n2290) );
  NAND2X1 U7227 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[15]), .B(en), 
        .Y(n2272) );
  OAI2BB1X1 U7228 ( 
        .A0N(output_p2_times_a2_div_componentxUDxquotient_not_gated[17]), 
        .A1N(n371), .B0(n2271), .Y(n2289) );
  NAND2X1 U7229 ( 
        .A(output_p2_times_a2_div_componentxUDxquotient_not_gated[16]), .B(en), 
        .Y(n2271) );
  INVX1 U7230 ( .A(n3570), .Y(n1451) );
  AOI22X1 U7231 ( .A0(input_p1_times_b1_div_componentxunsigned_output_11), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[11]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3570) );
  INVX1 U7232 ( .A(n3567), .Y(n1447) );
  AOI22X1 U7233 ( .A0(input_p1_times_b1_div_componentxunsigned_output_8), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[8]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3567) );
  INVX1 U7234 ( .A(n3561), .Y(n1441) );
  AOI22X1 U7235 ( .A0(input_p1_times_b1_div_componentxunsigned_output_2), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[2]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3561) );
  INVX1 U7236 ( .A(n3588), .Y(n1432) );
  AOI22X1 U7237 ( .A0(input_p2_times_b2_div_componentxunsigned_output_11), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[11]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3588) );
  INVX1 U7238 ( .A(n3585), .Y(n1428) );
  AOI22X1 U7239 ( .A0(input_p2_times_b2_div_componentxunsigned_output_8), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[8]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3585) );
  INVX1 U7240 ( .A(n3579), .Y(n1422) );
  AOI22X1 U7241 ( .A0(input_p2_times_b2_div_componentxunsigned_output_2), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[2]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3579) );
  INVX1 U7242 ( .A(n3606), .Y(n1413) );
  AOI22X1 U7243 ( .A0(output_p1_times_a1_div_componentxunsigned_output_11), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[11]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3606)
         );
  INVX1 U7244 ( .A(n3603), .Y(n1409) );
  AOI22X1 U7245 ( .A0(output_p1_times_a1_div_componentxunsigned_output_8), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[8]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3603)
         );
  INVX1 U7246 ( .A(n3597), .Y(n1403) );
  AOI22X1 U7247 ( .A0(output_p1_times_a1_div_componentxunsigned_output_2), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[2]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3597)
         );
  INVX1 U7248 ( .A(n3624), .Y(n1394) );
  AOI22X1 U7249 ( .A0(output_p2_times_a2_div_componentxunsigned_output_11), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[11]), 
        .B1(n7), .Y(n3624) );
  INVX1 U7250 ( .A(n3621), .Y(n1390) );
  AOI22X1 U7251 ( .A0(output_p2_times_a2_div_componentxunsigned_output_8), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[8]), 
        .B1(n7), .Y(n3621) );
  INVX1 U7252 ( .A(n3615), .Y(n1384) );
  AOI22X1 U7253 ( .A0(output_p2_times_a2_div_componentxunsigned_output_2), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[2]), 
        .B1(n7), .Y(n3615) );
  INVX1 U7254 ( .A(input_times_b0_div_componentxUDxn13), .Y(n1275) );
  AOI22X1 U7255 ( .A0(input_times_b0_div_componentxunsigned_output_11), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[11]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn13) );
  INVX1 U7256 ( .A(input_times_b0_div_componentxUDxn10), .Y(n1271) );
  AOI22X1 U7257 ( .A0(input_times_b0_div_componentxunsigned_output_8), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[8]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn10) );
  INVX1 U7258 ( .A(input_times_b0_div_componentxUDxn4), .Y(n1265) );
  AOI22X1 U7259 ( .A0(input_times_b0_div_componentxunsigned_output_2), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[2]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn4) );
  INVX1 U7260 ( .A(n3576), .Y(n1457) );
  AOI22X1 U7261 ( .A0(input_p1_times_b1_div_componentxunsigned_output_17), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[17]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3576) );
  INVX1 U7262 ( .A(n3575), .Y(n1456) );
  AOI22X1 U7263 ( .A0(input_p1_times_b1_div_componentxunsigned_output_16), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[16]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3575) );
  INVX1 U7264 ( .A(n3573), .Y(n1454) );
  AOI22X1 U7265 ( .A0(input_p1_times_b1_div_componentxunsigned_output_14), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[14]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3573) );
  INVX1 U7266 ( .A(n3572), .Y(n1453) );
  AOI22X1 U7267 ( .A0(input_p1_times_b1_div_componentxunsigned_output_13), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[13]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3572) );
  INVX1 U7268 ( .A(n3571), .Y(n1452) );
  AOI22X1 U7269 ( .A0(input_p1_times_b1_div_componentxunsigned_output_12), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[12]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3571) );
  INVX1 U7270 ( .A(n3569), .Y(n1450) );
  AOI22X1 U7271 ( .A0(input_p1_times_b1_div_componentxunsigned_output_10), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[10]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3569) );
  INVX1 U7272 ( .A(n3566), .Y(n1446) );
  AOI22X1 U7273 ( .A0(input_p1_times_b1_div_componentxunsigned_output_7), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[7]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3566) );
  INVX1 U7274 ( .A(n3564), .Y(n1444) );
  AOI22X1 U7275 ( .A0(input_p1_times_b1_div_componentxunsigned_output_5), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[5]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3564) );
  INVX1 U7276 ( .A(n3563), .Y(n1443) );
  AOI22X1 U7277 ( .A0(input_p1_times_b1_div_componentxunsigned_output_4), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[4]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3563) );
  INVX1 U7278 ( .A(n3562), .Y(n1442) );
  AOI22X1 U7279 ( .A0(input_p1_times_b1_div_componentxunsigned_output_3), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[3]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3562) );
  INVX1 U7280 ( .A(n3560), .Y(n1440) );
  AOI22X1 U7281 ( .A0(input_p1_times_b1_div_componentxunsigned_output_1), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[1]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3560) );
  INVX1 U7282 ( .A(n3559), .Y(n1439) );
  AOI22X1 U7283 ( 
        .A0(input_p1_times_b1_div_componentxunsigned_output_inverted[0]), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[0]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3559) );
  INVX1 U7284 ( .A(n3594), .Y(n1438) );
  AOI22X1 U7285 ( .A0(input_p2_times_b2_div_componentxunsigned_output_17), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[17]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3594) );
  INVX1 U7286 ( .A(n3593), .Y(n1437) );
  AOI22X1 U7287 ( .A0(input_p2_times_b2_div_componentxunsigned_output_16), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[16]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3593) );
  INVX1 U7288 ( .A(n3591), .Y(n1435) );
  AOI22X1 U7289 ( .A0(input_p2_times_b2_div_componentxunsigned_output_14), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[14]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3591) );
  INVX1 U7290 ( .A(n3590), .Y(n1434) );
  AOI22X1 U7291 ( .A0(input_p2_times_b2_div_componentxunsigned_output_13), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[13]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3590) );
  INVX1 U7292 ( .A(n3589), .Y(n1433) );
  AOI22X1 U7293 ( .A0(input_p2_times_b2_div_componentxunsigned_output_12), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[12]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3589) );
  INVX1 U7294 ( .A(n3587), .Y(n1431) );
  AOI22X1 U7295 ( .A0(input_p2_times_b2_div_componentxunsigned_output_10), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[10]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3587) );
  INVX1 U7296 ( .A(n3584), .Y(n1427) );
  AOI22X1 U7297 ( .A0(input_p2_times_b2_div_componentxunsigned_output_7), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[7]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3584) );
  INVX1 U7298 ( .A(n3582), .Y(n1425) );
  AOI22X1 U7299 ( .A0(input_p2_times_b2_div_componentxunsigned_output_5), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[5]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3582) );
  INVX1 U7300 ( .A(n3581), .Y(n1424) );
  AOI22X1 U7301 ( .A0(input_p2_times_b2_div_componentxunsigned_output_4), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[4]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3581) );
  INVX1 U7302 ( .A(n3580), .Y(n1423) );
  AOI22X1 U7303 ( .A0(input_p2_times_b2_div_componentxunsigned_output_3), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[3]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3580) );
  INVX1 U7304 ( .A(n3578), .Y(n1421) );
  AOI22X1 U7305 ( .A0(input_p2_times_b2_div_componentxunsigned_output_1), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[1]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3578) );
  INVX1 U7306 ( .A(n3577), .Y(n1420) );
  AOI22X1 U7307 ( 
        .A0(input_p2_times_b2_div_componentxunsigned_output_inverted[0]), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[0]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3577) );
  INVX1 U7308 ( .A(n3612), .Y(n1419) );
  AOI22X1 U7309 ( .A0(output_p1_times_a1_div_componentxunsigned_output_17), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[17]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3612)
         );
  INVX1 U7310 ( .A(n3611), .Y(n1418) );
  AOI22X1 U7311 ( .A0(output_p1_times_a1_div_componentxunsigned_output_16), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[16]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3611)
         );
  INVX1 U7312 ( .A(n3609), .Y(n1416) );
  AOI22X1 U7313 ( .A0(output_p1_times_a1_div_componentxunsigned_output_14), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[14]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3609)
         );
  INVX1 U7314 ( .A(n3608), .Y(n1415) );
  AOI22X1 U7315 ( .A0(output_p1_times_a1_div_componentxunsigned_output_13), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[13]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3608)
         );
  INVX1 U7316 ( .A(n3607), .Y(n1414) );
  AOI22X1 U7317 ( .A0(output_p1_times_a1_div_componentxunsigned_output_12), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[12]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3607)
         );
  INVX1 U7318 ( .A(n3605), .Y(n1412) );
  AOI22X1 U7319 ( .A0(output_p1_times_a1_div_componentxunsigned_output_10), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[10]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3605)
         );
  INVX1 U7320 ( .A(n3602), .Y(n1408) );
  AOI22X1 U7321 ( .A0(output_p1_times_a1_div_componentxunsigned_output_7), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[7]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3602)
         );
  INVX1 U7322 ( .A(n3600), .Y(n1406) );
  AOI22X1 U7323 ( .A0(output_p1_times_a1_div_componentxunsigned_output_5), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[5]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3600)
         );
  INVX1 U7324 ( .A(n3599), .Y(n1405) );
  AOI22X1 U7325 ( .A0(output_p1_times_a1_div_componentxunsigned_output_4), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[4]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3599)
         );
  INVX1 U7326 ( .A(n3598), .Y(n1404) );
  AOI22X1 U7327 ( .A0(output_p1_times_a1_div_componentxunsigned_output_3), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[3]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3598)
         );
  INVX1 U7328 ( .A(n3596), .Y(n1402) );
  AOI22X1 U7329 ( .A0(output_p1_times_a1_div_componentxunsigned_output_1), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[1]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3596)
         );
  INVX1 U7330 ( .A(n3595), .Y(n1401) );
  AOI22X1 U7331 ( 
        .A0(output_p1_times_a1_div_componentxunsigned_output_inverted[0]), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[0]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3595)
         );
  INVX1 U7332 ( .A(n3630), .Y(n1400) );
  AOI22X1 U7333 ( .A0(output_p2_times_a2_div_componentxunsigned_output_17), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[17]), 
        .B1(n7), .Y(n3630) );
  INVX1 U7334 ( .A(n3629), .Y(n1399) );
  AOI22X1 U7335 ( .A0(output_p2_times_a2_div_componentxunsigned_output_16), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[16]), 
        .B1(n7), .Y(n3629) );
  INVX1 U7336 ( .A(n3627), .Y(n1397) );
  AOI22X1 U7337 ( .A0(output_p2_times_a2_div_componentxunsigned_output_14), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[14]), 
        .B1(n7), .Y(n3627) );
  INVX1 U7338 ( .A(n3626), .Y(n1396) );
  AOI22X1 U7339 ( .A0(output_p2_times_a2_div_componentxunsigned_output_13), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[13]), 
        .B1(n7), .Y(n3626) );
  INVX1 U7340 ( .A(n3625), .Y(n1395) );
  AOI22X1 U7341 ( .A0(output_p2_times_a2_div_componentxunsigned_output_12), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[12]), 
        .B1(n7), .Y(n3625) );
  INVX1 U7342 ( .A(n3623), .Y(n1393) );
  AOI22X1 U7343 ( .A0(output_p2_times_a2_div_componentxunsigned_output_10), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[10]), 
        .B1(n7), .Y(n3623) );
  INVX1 U7344 ( .A(n3620), .Y(n1389) );
  AOI22X1 U7345 ( .A0(output_p2_times_a2_div_componentxunsigned_output_7), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[7]), 
        .B1(n7), .Y(n3620) );
  INVX1 U7346 ( .A(n3618), .Y(n1387) );
  AOI22X1 U7347 ( .A0(output_p2_times_a2_div_componentxunsigned_output_5), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[5]), 
        .B1(n7), .Y(n3618) );
  INVX1 U7348 ( .A(n3617), .Y(n1386) );
  AOI22X1 U7349 ( .A0(output_p2_times_a2_div_componentxunsigned_output_4), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[4]), 
        .B1(n7), .Y(n3617) );
  INVX1 U7350 ( .A(n3616), .Y(n1385) );
  AOI22X1 U7351 ( .A0(output_p2_times_a2_div_componentxunsigned_output_3), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[3]), 
        .B1(n7), .Y(n3616) );
  INVX1 U7352 ( .A(n3614), .Y(n1383) );
  AOI22X1 U7353 ( .A0(output_p2_times_a2_div_componentxunsigned_output_1), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[1]), 
        .B1(n7), .Y(n3614) );
  INVX1 U7354 ( .A(n3613), .Y(n1382) );
  AOI22X1 U7355 ( 
        .A0(output_p2_times_a2_div_componentxunsigned_output_inverted[0]), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[0]), 
        .B1(n7), .Y(n3613) );
  INVX1 U7356 ( .A(input_times_b0_div_componentxUDxn19), .Y(n1281) );
  AOI22X1 U7357 ( .A0(input_times_b0_div_componentxunsigned_output_17), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[17]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn19) );
  INVX1 U7358 ( .A(input_times_b0_div_componentxUDxn18), .Y(n1280) );
  AOI22X1 U7359 ( .A0(input_times_b0_div_componentxunsigned_output_16), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[16]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn18) );
  INVX1 U7360 ( .A(input_times_b0_div_componentxUDxn16), .Y(n1278) );
  AOI22X1 U7361 ( .A0(input_times_b0_div_componentxunsigned_output_14), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[14]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn16) );
  INVX1 U7362 ( .A(input_times_b0_div_componentxUDxn15), .Y(n1277) );
  AOI22X1 U7363 ( .A0(input_times_b0_div_componentxunsigned_output_13), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[13]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn15) );
  INVX1 U7364 ( .A(input_times_b0_div_componentxUDxn14), .Y(n1276) );
  AOI22X1 U7365 ( .A0(input_times_b0_div_componentxunsigned_output_12), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[12]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn14) );
  INVX1 U7366 ( .A(input_times_b0_div_componentxUDxn12), .Y(n1274) );
  AOI22X1 U7367 ( .A0(input_times_b0_div_componentxunsigned_output_10), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[10]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn12) );
  INVX1 U7368 ( .A(input_times_b0_div_componentxUDxn9), .Y(n1270) );
  AOI22X1 U7369 ( .A0(input_times_b0_div_componentxunsigned_output_7), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[7]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn9) );
  INVX1 U7370 ( .A(input_times_b0_div_componentxUDxn7), .Y(n1268) );
  AOI22X1 U7371 ( .A0(input_times_b0_div_componentxunsigned_output_5), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[5]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn7) );
  INVX1 U7372 ( .A(input_times_b0_div_componentxUDxn6), .Y(n1267) );
  AOI22X1 U7373 ( .A0(input_times_b0_div_componentxunsigned_output_4), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[4]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn6) );
  INVX1 U7374 ( .A(input_times_b0_div_componentxUDxn5), .Y(n1266) );
  AOI22X1 U7375 ( .A0(input_times_b0_div_componentxunsigned_output_3), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[3]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn5) );
  INVX1 U7376 ( .A(input_times_b0_div_componentxUDxn3), .Y(n1264) );
  AOI22X1 U7377 ( .A0(input_times_b0_div_componentxunsigned_output_1), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[1]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn3) );
  INVX1 U7378 ( .A(input_times_b0_div_componentxUDxn1), .Y(n1263) );
  AOI22X1 U7379 ( 
        .A0(input_times_b0_div_componentxunsigned_output_inverted[0]), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[0]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn1) );
  INVX1 U7380 ( .A(n3574), .Y(n1455) );
  AOI22X1 U7381 ( .A0(input_p1_times_b1_div_componentxunsigned_output_15), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[15]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3574) );
  INVX1 U7382 ( .A(n3568), .Y(n1449) );
  AOI22X1 U7383 ( .A0(input_p1_times_b1_div_componentxunsigned_output_9), 
        .A1(n159), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[9]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3568) );
  INVX1 U7384 ( .A(n3565), .Y(n1445) );
  AOI22X1 U7385 ( .A0(input_p1_times_b1_div_componentxunsigned_output_6), 
        .A1(n160), 
        .B0(input_p1_times_b1_div_componentxUDxquotient_not_gated[6]), 
        .B1(input_p1_times_b1_div_componentxoutput_ready_signal), .Y(n3565) );
  INVX1 U7386 ( .A(n3592), .Y(n1436) );
  AOI22X1 U7387 ( .A0(input_p2_times_b2_div_componentxunsigned_output_15), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[15]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3592) );
  INVX1 U7388 ( .A(n3586), .Y(n1430) );
  AOI22X1 U7389 ( .A0(input_p2_times_b2_div_componentxunsigned_output_9), 
        .A1(n157), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[9]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3586) );
  INVX1 U7390 ( .A(n3583), .Y(n1426) );
  AOI22X1 U7391 ( .A0(input_p2_times_b2_div_componentxunsigned_output_6), 
        .A1(n158), 
        .B0(input_p2_times_b2_div_componentxUDxquotient_not_gated[6]), 
        .B1(input_p2_times_b2_div_componentxoutput_ready_signal), .Y(n3583) );
  INVX1 U7392 ( .A(n3610), .Y(n1417) );
  AOI22X1 U7393 ( .A0(output_p1_times_a1_div_componentxunsigned_output_15), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[15]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3610)
         );
  INVX1 U7394 ( .A(n3604), .Y(n1411) );
  AOI22X1 U7395 ( .A0(output_p1_times_a1_div_componentxunsigned_output_9), 
        .A1(n155), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[9]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3604)
         );
  INVX1 U7396 ( .A(n3601), .Y(n1407) );
  AOI22X1 U7397 ( .A0(output_p1_times_a1_div_componentxunsigned_output_6), 
        .A1(n156), 
        .B0(output_p1_times_a1_div_componentxUDxquotient_not_gated[6]), 
        .B1(output_p1_times_a1_div_componentxoutput_ready_signal), .Y(n3601)
         );
  INVX1 U7398 ( .A(n3628), .Y(n1398) );
  AOI22X1 U7399 ( .A0(output_p2_times_a2_div_componentxunsigned_output_15), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[15]), 
        .B1(n7), .Y(n3628) );
  INVX1 U7400 ( .A(n3622), .Y(n1392) );
  AOI22X1 U7401 ( .A0(output_p2_times_a2_div_componentxunsigned_output_9), 
        .A1(n153), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[9]), 
        .B1(n7), .Y(n3622) );
  INVX1 U7402 ( .A(n3619), .Y(n1388) );
  AOI22X1 U7403 ( .A0(output_p2_times_a2_div_componentxunsigned_output_6), 
        .A1(n154), 
        .B0(output_p2_times_a2_div_componentxUDxquotient_not_gated[6]), 
        .B1(n7), .Y(n3619) );
  INVX1 U7404 ( .A(input_times_b0_div_componentxUDxn17), .Y(n1279) );
  AOI22X1 U7405 ( .A0(input_times_b0_div_componentxunsigned_output_15), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[15]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn17) );
  INVX1 U7406 ( .A(input_times_b0_div_componentxUDxn11), .Y(n1273) );
  AOI22X1 U7407 ( .A0(input_times_b0_div_componentxunsigned_output_9), 
        .A1(n137), .B0(input_times_b0_div_componentxUDxquotient_not_gated[9]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn11) );
  INVX1 U7408 ( .A(input_times_b0_div_componentxUDxn8), .Y(n1269) );
  AOI22X1 U7409 ( .A0(input_times_b0_div_componentxunsigned_output_6), 
        .A1(n138), .B0(input_times_b0_div_componentxUDxquotient_not_gated[6]), 
        .B1(n8), .Y(input_times_b0_div_componentxUDxn8) );
  AOI22X1 U7410 ( .A0(\parameter_B0_div[2] ), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_2_), .B1(n341), 
        .Y(input_times_b0_div_componentxn47) );
  XNOR2X1 U7411 ( .A(\parameter_B0_div[2] ), .B(n3889), 
        .Y(input_times_b0_div_componentxinput_B_inverted_2_) );
  NOR2X1 U7412 ( .A(\parameter_B0_div[0] ), .B(\parameter_B0_div[1] ), 
        .Y(n3889) );
  AOI22X1 U7413 ( .A0(\parameter_B1_div[2] ), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_2_), .B1(n332), 
        .Y(n4225) );
  XNOR2X1 U7414 ( .A(\parameter_B1_div[2] ), .B(n3932), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_2_) );
  NOR2X1 U7415 ( .A(\parameter_B1_div[0] ), .B(\parameter_B1_div[1] ), 
        .Y(n3932) );
  AOI22X1 U7416 ( .A0(\parameter_B2_div[2] ), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_2_), .B1(n323), 
        .Y(n4281) );
  XNOR2X1 U7417 ( .A(\parameter_B2_div[2] ), .B(n3975), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_2_) );
  NOR2X1 U7418 ( .A(\parameter_B2_div[0] ), .B(\parameter_B2_div[1] ), 
        .Y(n3975) );
  AOI22X1 U7419 ( .A0(\parameter_A1_div[2] ), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_2_), .B1(n359), 
        .Y(n4335) );
  XNOR2X1 U7420 ( .A(\parameter_A1_div[2] ), .B(n4018), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_2_) );
  NOR2X1 U7421 ( .A(\parameter_A1_div[0] ), .B(\parameter_A1_div[1] ), 
        .Y(n4018) );
  AOI22X1 U7422 ( .A0(\parameter_A2_div[2] ), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_2_), .B1(n350), 
        .Y(n4391) );
  XNOR2X1 U7423 ( .A(\parameter_A2_div[2] ), .B(n4061), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_2_) );
  NOR2X1 U7424 ( .A(\parameter_A2_div[0] ), .B(\parameter_A2_div[1] ), 
        .Y(n4061) );
  AOI22X1 U7425 ( .A0(\parameter_B0_div[4] ), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_4_), .B1(n341), 
        .Y(input_times_b0_div_componentxn49) );
  XOR2X1 U7426 ( .A(n3887), .B(\parameter_B0_div[4] ), 
        .Y(input_times_b0_div_componentxinput_B_inverted_4_) );
  OR2X2 U7427 ( .A(\parameter_B0_div[3] ), .B(n3888), .Y(n3887) );
  AOI22X1 U7428 ( .A0(\parameter_B1_div[4] ), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_4_), .B1(n332), 
        .Y(n4227) );
  XOR2X1 U7429 ( .A(n3930), .B(\parameter_B1_div[4] ), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_4_) );
  OR2X2 U7430 ( .A(\parameter_B1_div[3] ), .B(n3931), .Y(n3930) );
  AOI22X1 U7431 ( .A0(\parameter_B2_div[4] ), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_4_), .B1(n323), 
        .Y(n4283) );
  XOR2X1 U7432 ( .A(n3973), .B(\parameter_B2_div[4] ), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_4_) );
  OR2X2 U7433 ( .A(\parameter_B2_div[3] ), .B(n3974), .Y(n3973) );
  AOI22X1 U7434 ( .A0(\parameter_A1_div[4] ), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_4_), .B1(n359), 
        .Y(n4337) );
  XOR2X1 U7435 ( .A(n4016), .B(\parameter_A1_div[4] ), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_4_) );
  OR2X2 U7436 ( .A(\parameter_A1_div[3] ), .B(n4017), .Y(n4016) );
  AOI22X1 U7437 ( .A0(\parameter_A2_div[4] ), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_4_), .B1(n350), 
        .Y(n4393) );
  XOR2X1 U7438 ( .A(n4059), .B(\parameter_A2_div[4] ), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_4_) );
  OR2X2 U7439 ( .A(\parameter_A2_div[3] ), .B(n4060), .Y(n4059) );
  AOI22X1 U7440 ( .A0(\parameter_B0_div[6] ), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_6_), .B1(n341), 
        .Y(input_times_b0_div_componentxn51) );
  XOR2X1 U7441 ( .A(n3885), .B(\parameter_B0_div[6] ), 
        .Y(input_times_b0_div_componentxinput_B_inverted_6_) );
  OR2X2 U7442 ( .A(\parameter_B0_div[5] ), .B(n3886), .Y(n3885) );
  AOI22X1 U7443 ( .A0(\parameter_B1_div[6] ), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_6_), .B1(n332), 
        .Y(n4229) );
  XOR2X1 U7444 ( .A(n3928), .B(\parameter_B1_div[6] ), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_6_) );
  OR2X2 U7445 ( .A(\parameter_B1_div[5] ), .B(n3929), .Y(n3928) );
  AOI22X1 U7446 ( .A0(\parameter_B2_div[6] ), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_6_), .B1(n323), 
        .Y(n4285) );
  XOR2X1 U7447 ( .A(n3971), .B(\parameter_B2_div[6] ), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_6_) );
  OR2X2 U7448 ( .A(\parameter_B2_div[5] ), .B(n3972), .Y(n3971) );
  AOI22X1 U7449 ( .A0(\parameter_A1_div[6] ), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_6_), .B1(n359), 
        .Y(n4339) );
  XOR2X1 U7450 ( .A(n4014), .B(\parameter_A1_div[6] ), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_6_) );
  OR2X2 U7451 ( .A(\parameter_A1_div[5] ), .B(n4015), .Y(n4014) );
  AOI22X1 U7452 ( .A0(\parameter_A2_div[6] ), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_6_), .B1(n350), 
        .Y(n4395) );
  XOR2X1 U7453 ( .A(n4057), .B(\parameter_A2_div[6] ), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_6_) );
  OR2X2 U7454 ( .A(\parameter_A2_div[5] ), .B(n4058), .Y(n4057) );
  AOI22X1 U7455 ( .A0(\parameter_B0_div[3] ), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_3_), .B1(n341), 
        .Y(input_times_b0_div_componentxn48) );
  XOR2X1 U7456 ( .A(n3888), .B(\parameter_B0_div[3] ), 
        .Y(input_times_b0_div_componentxinput_B_inverted_3_) );
  AOI22X1 U7457 ( .A0(\parameter_B1_div[3] ), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_3_), .B1(n332), 
        .Y(n4226) );
  XOR2X1 U7458 ( .A(n3931), .B(\parameter_B1_div[3] ), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_3_) );
  AOI22X1 U7459 ( .A0(\parameter_B2_div[3] ), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_3_), .B1(n323), 
        .Y(n4282) );
  XOR2X1 U7460 ( .A(n3974), .B(\parameter_B2_div[3] ), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_3_) );
  AOI22X1 U7461 ( .A0(\parameter_A1_div[3] ), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_3_), .B1(n359), 
        .Y(n4336) );
  XOR2X1 U7462 ( .A(n4017), .B(\parameter_A1_div[3] ), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_3_) );
  AOI22X1 U7463 ( .A0(\parameter_A2_div[3] ), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_3_), .B1(n350), 
        .Y(n4392) );
  XOR2X1 U7464 ( .A(n4060), .B(\parameter_A2_div[3] ), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_3_) );
  AOI22X1 U7465 ( .A0(\parameter_B0_div[5] ), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_5_), .B1(n341), 
        .Y(input_times_b0_div_componentxn50) );
  XOR2X1 U7466 ( .A(n3886), .B(\parameter_B0_div[5] ), 
        .Y(input_times_b0_div_componentxinput_B_inverted_5_) );
  AOI22X1 U7467 ( .A0(\parameter_B1_div[5] ), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_5_), .B1(n332), 
        .Y(n4228) );
  XOR2X1 U7468 ( .A(n3929), .B(\parameter_B1_div[5] ), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_5_) );
  AOI22X1 U7469 ( .A0(\parameter_B2_div[5] ), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_5_), .B1(n323), 
        .Y(n4284) );
  XOR2X1 U7470 ( .A(n3972), .B(\parameter_B2_div[5] ), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_5_) );
  AOI22X1 U7471 ( .A0(\parameter_A1_div[5] ), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_5_), .B1(n359), 
        .Y(n4338) );
  XOR2X1 U7472 ( .A(n4015), .B(\parameter_A1_div[5] ), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_5_) );
  AOI22X1 U7473 ( .A0(\parameter_A2_div[5] ), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_5_), .B1(n350), 
        .Y(n4394) );
  XOR2X1 U7474 ( .A(n4058), .B(\parameter_A2_div[5] ), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_5_) );
  INVX1 U7475 ( .A(input_times_b0_div_componentxn45), .Y(n846) );
  AOI22X1 U7476 ( .A0(\parameter_B0_div[0] ), .A1(n342), 
        .B0(\parameter_B0_div[0] ), .B1(n341), 
        .Y(input_times_b0_div_componentxn45) );
  INVX1 U7477 ( .A(n4223), .Y(n1005) );
  AOI22X1 U7478 ( .A0(\parameter_B1_div[0] ), .A1(n333), 
        .B0(\parameter_B1_div[0] ), .B1(n332), .Y(n4223) );
  INVX1 U7479 ( .A(n4279), .Y(n1164) );
  AOI22X1 U7480 ( .A0(\parameter_B2_div[0] ), .A1(n324), 
        .B0(\parameter_B2_div[0] ), .B1(n323), .Y(n4279) );
  INVX1 U7481 ( .A(n4333), .Y(n528) );
  AOI22X1 U7482 ( .A0(\parameter_A1_div[0] ), .A1(n360), 
        .B0(\parameter_A1_div[0] ), .B1(n359), .Y(n4333) );
  INVX1 U7483 ( .A(n4389), .Y(n687) );
  AOI22X1 U7484 ( .A0(\parameter_A2_div[0] ), .A1(n351), 
        .B0(\parameter_A2_div[0] ), .B1(n350), .Y(n4389) );
  OR3XL U7485 ( .A(\parameter_B1_mul[5] ), .B(\parameter_B1_mul[6] ), 
        .C(n3699), .Y(n3697) );
  OR3XL U7486 ( .A(\parameter_B2_mul[5] ), .B(\parameter_B2_mul[6] ), 
        .C(n3747), .Y(n3745) );
  OR3XL U7487 ( .A(\parameter_A2_mul[5] ), .B(\parameter_A2_mul[6] ), 
        .C(n3843), .Y(n3841) );
  OR3XL U7488 ( .A(\parameter_B0_mul[5] ), .B(\parameter_B0_mul[6] ), 
        .C(n3651), .Y(n3649) );
  OR3XL U7489 ( .A(\parameter_A1_mul[5] ), .B(\parameter_A1_mul[6] ), 
        .C(n3795), .Y(n3793) );
  OR3XL U7490 ( .A(\parameter_B0_div[5] ), .B(\parameter_B0_div[6] ), 
        .C(n3886), .Y(n3884) );
  OR3XL U7491 ( .A(\parameter_B1_div[5] ), .B(\parameter_B1_div[6] ), 
        .C(n3929), .Y(n3927) );
  OR3XL U7492 ( .A(\parameter_B2_div[5] ), .B(\parameter_B2_div[6] ), 
        .C(n3972), .Y(n3970) );
  OR3XL U7493 ( .A(\parameter_A1_div[5] ), .B(\parameter_A1_div[6] ), 
        .C(n4015), .Y(n4013) );
  OR3XL U7494 ( .A(\parameter_A2_div[5] ), .B(\parameter_A2_div[6] ), 
        .C(n4058), .Y(n4056) );
  OR3XL U7495 ( .A(\parameter_B1_mul[3] ), .B(\parameter_B1_mul[4] ), 
        .C(n3701), .Y(n3699) );
  OR3XL U7496 ( .A(\parameter_B2_mul[3] ), .B(\parameter_B2_mul[4] ), 
        .C(n3749), .Y(n3747) );
  OR3XL U7497 ( .A(\parameter_A2_mul[3] ), .B(\parameter_A2_mul[4] ), 
        .C(n3845), .Y(n3843) );
  OR3XL U7498 ( .A(\parameter_B0_mul[3] ), .B(\parameter_B0_mul[4] ), 
        .C(n3653), .Y(n3651) );
  OR3XL U7499 ( .A(\parameter_B0_div[3] ), .B(\parameter_B0_div[4] ), 
        .C(n3888), .Y(n3886) );
  OR3XL U7500 ( .A(\parameter_B1_div[3] ), .B(\parameter_B1_div[4] ), 
        .C(n3931), .Y(n3929) );
  OR3XL U7501 ( .A(\parameter_B2_div[3] ), .B(\parameter_B2_div[4] ), 
        .C(n3974), .Y(n3972) );
  OR3XL U7502 ( .A(\parameter_A1_mul[3] ), .B(\parameter_A1_mul[4] ), 
        .C(n3797), .Y(n3795) );
  OR3XL U7503 ( .A(\parameter_A1_div[3] ), .B(\parameter_A1_div[4] ), 
        .C(n4017), .Y(n4015) );
  OR3XL U7504 ( .A(\parameter_A2_div[3] ), .B(\parameter_A2_div[4] ), 
        .C(n4060), .Y(n4058) );
  OR3XL U7505 ( .A(\parameter_B1_mul[1] ), .B(\parameter_B1_mul[2] ), 
        .C(\parameter_B1_mul[0] ), .Y(n3701) );
  OR3XL U7506 ( .A(\parameter_B2_mul[1] ), .B(\parameter_B2_mul[2] ), 
        .C(\parameter_B2_mul[0] ), .Y(n3749) );
  OR3XL U7507 ( .A(\parameter_A1_mul[1] ), .B(\parameter_A1_mul[2] ), 
        .C(\parameter_A1_mul[0] ), .Y(n3797) );
  OR3XL U7508 ( .A(\parameter_A2_mul[1] ), .B(\parameter_A2_mul[2] ), 
        .C(\parameter_A2_mul[0] ), .Y(n3845) );
  OR3XL U7509 ( .A(\parameter_B0_mul[1] ), .B(\parameter_B0_mul[2] ), 
        .C(\parameter_B0_mul[0] ), .Y(n3653) );
  OR3XL U7510 ( .A(\parameter_B0_div[1] ), .B(\parameter_B0_div[2] ), 
        .C(\parameter_B0_div[0] ), .Y(n3888) );
  OR3XL U7511 ( .A(\parameter_B1_div[1] ), .B(\parameter_B1_div[2] ), 
        .C(\parameter_B1_div[0] ), .Y(n3931) );
  OR3XL U7512 ( .A(\parameter_B2_div[1] ), .B(\parameter_B2_div[2] ), 
        .C(\parameter_B2_div[0] ), .Y(n3974) );
  OR3XL U7513 ( .A(\parameter_A1_div[1] ), .B(\parameter_A1_div[2] ), 
        .C(\parameter_A1_div[0] ), .Y(n4017) );
  OR3XL U7514 ( .A(\parameter_A2_div[1] ), .B(\parameter_A2_div[2] ), 
        .C(\parameter_A2_div[0] ), .Y(n4060) );
  BUFX3 U7515 ( .A(n4423), .Y(n179) );
  AOI22X1 U7516 ( .A0(\parameter_B1_mul[0] ), .A1(n339), 
        .B0(\parameter_B1_mul[0] ), .B1(n336), .Y(n4423) );
  BUFX3 U7517 ( .A(n4476), .Y(n200) );
  AOI22X1 U7518 ( .A0(\parameter_B2_mul[0] ), .A1(n330), 
        .B0(\parameter_B2_mul[0] ), .B1(n327), .Y(n4476) );
  BUFX3 U7519 ( .A(n4582), .Y(n242) );
  AOI22X1 U7520 ( .A0(\parameter_A2_mul[0] ), .A1(n357), 
        .B0(\parameter_A2_mul[0] ), .B1(n354), .Y(n4582) );
  BUFX3 U7521 ( .A(input_times_b0_mul_componentxn72), .Y(n270) );
  AOI22X1 U7522 ( .A0(\parameter_B0_mul[0] ), .A1(n348), 
        .B0(\parameter_B0_mul[0] ), .B1(n345), 
        .Y(input_times_b0_mul_componentxn72) );
  BUFX3 U7523 ( .A(n4529), .Y(n221) );
  AOI22X1 U7524 ( .A0(\parameter_A1_mul[0] ), .A1(n366), 
        .B0(\parameter_A1_mul[0] ), .B1(n363), .Y(n4529) );
  BUFX3 U7525 ( .A(n4415), .Y(n178) );
  AOI22X1 U7526 ( .A0(\parameter_B1_mul[1] ), .A1(n338), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_1_), .B1(n335), 
        .Y(n4415) );
  XOR2X1 U7527 ( .A(\parameter_B1_mul[1] ), .B(\parameter_B1_mul[0] ), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_1_) );
  BUFX3 U7528 ( .A(n4468), .Y(n199) );
  AOI22X1 U7529 ( .A0(\parameter_B2_mul[1] ), .A1(n329), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_1_), .B1(n326), 
        .Y(n4468) );
  XOR2X1 U7530 ( .A(\parameter_B2_mul[1] ), .B(\parameter_B2_mul[0] ), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_1_) );
  BUFX3 U7531 ( .A(n4521), .Y(n220) );
  AOI22X1 U7532 ( .A0(\parameter_A1_mul[1] ), .A1(n365), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_1_), .B1(n362), 
        .Y(n4521) );
  XOR2X1 U7533 ( .A(\parameter_A1_mul[1] ), .B(\parameter_A1_mul[0] ), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_1_) );
  BUFX3 U7534 ( .A(n4574), .Y(n241) );
  AOI22X1 U7535 ( .A0(\parameter_A2_mul[1] ), .A1(n356), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_1_), .B1(n353), 
        .Y(n4574) );
  XOR2X1 U7536 ( .A(\parameter_A2_mul[1] ), .B(\parameter_A2_mul[0] ), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_1_) );
  BUFX3 U7537 ( .A(input_times_b0_mul_componentxn64), .Y(n269) );
  AOI22X1 U7538 ( .A0(\parameter_B0_mul[1] ), .A1(n347), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_1_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn64) );
  XOR2X1 U7539 ( .A(\parameter_B0_mul[1] ), .B(\parameter_B0_mul[0] ), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_1_) );
  BUFX3 U7540 ( .A(n4414), .Y(n177) );
  AOI22X1 U7541 ( .A0(\parameter_B1_mul[2] ), .A1(n338), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_2_), .B1(n335), 
        .Y(n4414) );
  XNOR2X1 U7542 ( .A(\parameter_B1_mul[2] ), .B(n3702), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_2_) );
  NOR2X1 U7543 ( .A(\parameter_B1_mul[0] ), .B(\parameter_B1_mul[1] ), 
        .Y(n3702) );
  BUFX3 U7544 ( .A(n4467), .Y(n198) );
  AOI22X1 U7545 ( .A0(\parameter_B2_mul[2] ), .A1(n329), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_2_), .B1(n326), 
        .Y(n4467) );
  XNOR2X1 U7546 ( .A(\parameter_B2_mul[2] ), .B(n3750), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_2_) );
  NOR2X1 U7547 ( .A(\parameter_B2_mul[0] ), .B(\parameter_B2_mul[1] ), 
        .Y(n3750) );
  BUFX3 U7548 ( .A(n4520), .Y(n219) );
  AOI22X1 U7549 ( .A0(\parameter_A1_mul[2] ), .A1(n365), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_2_), .B1(n362), 
        .Y(n4520) );
  XNOR2X1 U7550 ( .A(\parameter_A1_mul[2] ), .B(n3798), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_2_) );
  NOR2X1 U7551 ( .A(\parameter_A1_mul[0] ), .B(\parameter_A1_mul[1] ), 
        .Y(n3798) );
  BUFX3 U7552 ( .A(n4573), .Y(n240) );
  AOI22X1 U7553 ( .A0(\parameter_A2_mul[2] ), .A1(n356), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_2_), .B1(n353), 
        .Y(n4573) );
  XNOR2X1 U7554 ( .A(\parameter_A2_mul[2] ), .B(n3846), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_2_) );
  NOR2X1 U7555 ( .A(\parameter_A2_mul[0] ), .B(\parameter_A2_mul[1] ), 
        .Y(n3846) );
  BUFX3 U7556 ( .A(input_times_b0_mul_componentxn63), .Y(n268) );
  AOI22X1 U7557 ( .A0(\parameter_B0_mul[2] ), .A1(n347), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_2_), .B1(n345), 
        .Y(input_times_b0_mul_componentxn63) );
  XNOR2X1 U7558 ( .A(\parameter_B0_mul[2] ), .B(n3654), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_2_) );
  NOR2X1 U7559 ( .A(\parameter_B0_mul[0] ), .B(\parameter_B0_mul[1] ), 
        .Y(n3654) );
  BUFX3 U7560 ( .A(n4413), .Y(n176) );
  AOI22X1 U7561 ( .A0(\parameter_B1_mul[3] ), .A1(n339), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_3_), .B1(n335), 
        .Y(n4413) );
  XOR2X1 U7562 ( .A(n3701), .B(\parameter_B1_mul[3] ), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_3_) );
  BUFX3 U7563 ( .A(n4466), .Y(n197) );
  AOI22X1 U7564 ( .A0(\parameter_B2_mul[3] ), .A1(n330), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_3_), .B1(n326), 
        .Y(n4466) );
  XOR2X1 U7565 ( .A(n3749), .B(\parameter_B2_mul[3] ), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_3_) );
  BUFX3 U7566 ( .A(n4519), .Y(n218) );
  AOI22X1 U7567 ( .A0(\parameter_A1_mul[3] ), .A1(n366), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_3_), .B1(n362), 
        .Y(n4519) );
  XOR2X1 U7568 ( .A(n3797), .B(\parameter_A1_mul[3] ), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_3_) );
  BUFX3 U7569 ( .A(n4572), .Y(n239) );
  AOI22X1 U7570 ( .A0(\parameter_A2_mul[3] ), .A1(n357), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_3_), .B1(n353), 
        .Y(n4572) );
  XOR2X1 U7571 ( .A(n3845), .B(\parameter_A2_mul[3] ), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_3_) );
  BUFX3 U7572 ( .A(input_times_b0_mul_componentxn62), .Y(n267) );
  AOI22X1 U7573 ( .A0(\parameter_B0_mul[3] ), .A1(n348), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_3_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn62) );
  XOR2X1 U7574 ( .A(n3653), .B(\parameter_B0_mul[3] ), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_3_) );
  INVX1 U7575 ( .A(en), .Y(n368) );
  BUFX3 U7576 ( .A(n4412), .Y(n175) );
  AOI22X1 U7577 ( .A0(\parameter_B1_mul[4] ), .A1(n338), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_4_), .B1(n335), 
        .Y(n4412) );
  XOR2X1 U7578 ( .A(n3700), .B(\parameter_B1_mul[4] ), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_4_) );
  OR2X2 U7579 ( .A(\parameter_B1_mul[3] ), .B(n3701), .Y(n3700) );
  BUFX3 U7580 ( .A(n4465), .Y(n196) );
  AOI22X1 U7581 ( .A0(\parameter_B2_mul[4] ), .A1(n329), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_4_), .B1(n326), 
        .Y(n4465) );
  XOR2X1 U7582 ( .A(n3748), .B(\parameter_B2_mul[4] ), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_4_) );
  OR2X2 U7583 ( .A(\parameter_B2_mul[3] ), .B(n3749), .Y(n3748) );
  BUFX3 U7584 ( .A(n4518), .Y(n217) );
  AOI22X1 U7585 ( .A0(\parameter_A1_mul[4] ), .A1(n365), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_4_), .B1(n362), 
        .Y(n4518) );
  XOR2X1 U7586 ( .A(n3796), .B(\parameter_A1_mul[4] ), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_4_) );
  OR2X2 U7587 ( .A(\parameter_A1_mul[3] ), .B(n3797), .Y(n3796) );
  BUFX3 U7588 ( .A(n4571), .Y(n238) );
  AOI22X1 U7589 ( .A0(\parameter_A2_mul[4] ), .A1(n356), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_4_), .B1(n353), 
        .Y(n4571) );
  XOR2X1 U7590 ( .A(n3844), .B(\parameter_A2_mul[4] ), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_4_) );
  OR2X2 U7591 ( .A(\parameter_A2_mul[3] ), .B(n3845), .Y(n3844) );
  BUFX3 U7592 ( .A(input_times_b0_mul_componentxn61), .Y(n266) );
  AOI22X1 U7593 ( .A0(\parameter_B0_mul[4] ), .A1(n347), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_4_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn61) );
  XOR2X1 U7594 ( .A(n3652), .B(\parameter_B0_mul[4] ), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_4_) );
  OR2X2 U7595 ( .A(\parameter_B0_mul[3] ), .B(n3653), .Y(n3652) );
  INVX1 U7596 ( .A(input_times_b0_div_componentxn46), .Y(n847) );
  AOI22X1 U7597 ( .A0(\parameter_B0_div[1] ), .A1(n342), 
        .B0(input_times_b0_div_componentxinput_B_inverted_1_), .B1(n341), 
        .Y(input_times_b0_div_componentxn46) );
  XOR2X1 U7598 ( .A(\parameter_B0_div[1] ), .B(\parameter_B0_div[0] ), 
        .Y(input_times_b0_div_componentxinput_B_inverted_1_) );
  INVX1 U7599 ( .A(n4224), .Y(n1006) );
  AOI22X1 U7600 ( .A0(\parameter_B1_div[1] ), .A1(n333), 
        .B0(input_p1_times_b1_div_componentxinput_B_inverted_1_), .B1(n332), 
        .Y(n4224) );
  XOR2X1 U7601 ( .A(\parameter_B1_div[1] ), .B(\parameter_B1_div[0] ), 
        .Y(input_p1_times_b1_div_componentxinput_B_inverted_1_) );
  INVX1 U7602 ( .A(n4280), .Y(n1165) );
  AOI22X1 U7603 ( .A0(\parameter_B2_div[1] ), .A1(n324), 
        .B0(input_p2_times_b2_div_componentxinput_B_inverted_1_), .B1(n323), 
        .Y(n4280) );
  XOR2X1 U7604 ( .A(\parameter_B2_div[1] ), .B(\parameter_B2_div[0] ), 
        .Y(input_p2_times_b2_div_componentxinput_B_inverted_1_) );
  INVX1 U7605 ( .A(n4334), .Y(n529) );
  AOI22X1 U7606 ( .A0(\parameter_A1_div[1] ), .A1(n360), 
        .B0(output_p1_times_a1_div_componentxinput_B_inverted_1_), .B1(n359), 
        .Y(n4334) );
  XOR2X1 U7607 ( .A(\parameter_A1_div[1] ), .B(\parameter_A1_div[0] ), 
        .Y(output_p1_times_a1_div_componentxinput_B_inverted_1_) );
  INVX1 U7608 ( .A(n4390), .Y(n688) );
  AOI22X1 U7609 ( .A0(\parameter_A2_div[1] ), .A1(n351), 
        .B0(output_p2_times_a2_div_componentxinput_B_inverted_1_), .B1(n350), 
        .Y(n4390) );
  XOR2X1 U7610 ( .A(\parameter_A2_div[1] ), .B(\parameter_A2_div[0] ), 
        .Y(output_p2_times_a2_div_componentxinput_B_inverted_1_) );
  BUFX3 U7611 ( .A(n4411), .Y(n174) );
  AOI22X1 U7612 ( .A0(\parameter_B1_mul[5] ), .A1(n339), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_5_), .B1(n335), 
        .Y(n4411) );
  XOR2X1 U7613 ( .A(n3699), .B(\parameter_B1_mul[5] ), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_5_) );
  BUFX3 U7614 ( .A(n4464), .Y(n195) );
  AOI22X1 U7615 ( .A0(\parameter_B2_mul[5] ), .A1(n330), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_5_), .B1(n326), 
        .Y(n4464) );
  XOR2X1 U7616 ( .A(n3747), .B(\parameter_B2_mul[5] ), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_5_) );
  BUFX3 U7617 ( .A(n4517), .Y(n216) );
  AOI22X1 U7618 ( .A0(\parameter_A1_mul[5] ), .A1(n366), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_5_), .B1(n362), 
        .Y(n4517) );
  XOR2X1 U7619 ( .A(n3795), .B(\parameter_A1_mul[5] ), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_5_) );
  BUFX3 U7620 ( .A(n4570), .Y(n237) );
  AOI22X1 U7621 ( .A0(\parameter_A2_mul[5] ), .A1(n357), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_5_), .B1(n353), 
        .Y(n4570) );
  XOR2X1 U7622 ( .A(n3843), .B(\parameter_A2_mul[5] ), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_5_) );
  BUFX3 U7623 ( .A(input_times_b0_mul_componentxn60), .Y(n265) );
  AOI22X1 U7624 ( .A0(\parameter_B0_mul[5] ), .A1(n348), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_5_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn60) );
  XOR2X1 U7625 ( .A(n3651), .B(\parameter_B0_mul[5] ), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_5_) );
  INVX1 U7626 ( .A(n337), .Y(n336) );
  INVX1 U7627 ( .A(n328), .Y(n327) );
  INVX1 U7628 ( .A(n355), .Y(n354) );
  INVX1 U7629 ( .A(n346), .Y(n345) );
  INVX1 U7630 ( .A(n364), .Y(n363) );
  BUFX3 U7631 ( .A(n4410), .Y(n173) );
  AOI22X1 U7632 ( .A0(\parameter_B1_mul[6] ), .A1(n338), 
        .B0(input_p1_times_b1_mul_componentxinput_B_inverted_6_), .B1(n335), 
        .Y(n4410) );
  XOR2X1 U7633 ( .A(n3698), .B(\parameter_B1_mul[6] ), 
        .Y(input_p1_times_b1_mul_componentxinput_B_inverted_6_) );
  OR2X2 U7634 ( .A(\parameter_B1_mul[5] ), .B(n3699), .Y(n3698) );
  BUFX3 U7635 ( .A(n4463), .Y(n194) );
  AOI22X1 U7636 ( .A0(\parameter_B2_mul[6] ), .A1(n329), 
        .B0(input_p2_times_b2_mul_componentxinput_B_inverted_6_), .B1(n326), 
        .Y(n4463) );
  XOR2X1 U7637 ( .A(n3746), .B(\parameter_B2_mul[6] ), 
        .Y(input_p2_times_b2_mul_componentxinput_B_inverted_6_) );
  OR2X2 U7638 ( .A(\parameter_B2_mul[5] ), .B(n3747), .Y(n3746) );
  BUFX3 U7639 ( .A(n4516), .Y(n215) );
  AOI22X1 U7640 ( .A0(\parameter_A1_mul[6] ), .A1(n365), 
        .B0(output_p1_times_a1_mul_componentxinput_B_inverted_6_), .B1(n362), 
        .Y(n4516) );
  XOR2X1 U7641 ( .A(n3794), .B(\parameter_A1_mul[6] ), 
        .Y(output_p1_times_a1_mul_componentxinput_B_inverted_6_) );
  OR2X2 U7642 ( .A(\parameter_A1_mul[5] ), .B(n3795), .Y(n3794) );
  BUFX3 U7643 ( .A(n4569), .Y(n236) );
  AOI22X1 U7644 ( .A0(\parameter_A2_mul[6] ), .A1(n356), 
        .B0(output_p2_times_a2_mul_componentxinput_B_inverted_6_), .B1(n353), 
        .Y(n4569) );
  XOR2X1 U7645 ( .A(n3842), .B(\parameter_A2_mul[6] ), 
        .Y(output_p2_times_a2_mul_componentxinput_B_inverted_6_) );
  OR2X2 U7646 ( .A(\parameter_A2_mul[5] ), .B(n3843), .Y(n3842) );
  BUFX3 U7647 ( .A(input_times_b0_mul_componentxn59), .Y(n264) );
  AOI22X1 U7648 ( .A0(\parameter_B0_mul[6] ), .A1(n347), 
        .B0(input_times_b0_mul_componentxinput_B_inverted_6_), .B1(n344), 
        .Y(input_times_b0_mul_componentxn59) );
  XOR2X1 U7649 ( .A(n3650), .B(\parameter_B0_mul[6] ), 
        .Y(input_times_b0_mul_componentxinput_B_inverted_6_) );
  OR2X2 U7650 ( .A(\parameter_B0_mul[5] ), .B(n3651), .Y(n3650) );
  INVX1 U7651 ( .A(\input_signal[7] ), .Y(n1174) );
  INVX1 U7652 ( .A(\parameter_B0_div[7] ), .Y(n342) );
  INVX1 U7653 ( .A(\parameter_B1_div[7] ), .Y(n333) );
  INVX1 U7654 ( .A(\parameter_B2_div[7] ), .Y(n324) );
  INVX1 U7655 ( .A(\parameter_A1_div[7] ), .Y(n360) );
  INVX1 U7656 ( .A(\parameter_A2_div[7] ), .Y(n351) );
  INVX1 U7657 ( .A(\parameter_B1_mul[7] ), .Y(n339) );
  INVX1 U7658 ( .A(\parameter_B2_mul[7] ), .Y(n330) );
  INVX1 U7659 ( .A(\parameter_A2_mul[7] ), .Y(n357) );
  INVX1 U7660 ( .A(\parameter_A1_mul[7] ), .Y(n366) );
  INVX1 U7661 ( .A(\parameter_B0_mul[7] ), .Y(n348) );
  INVX1 U7662 ( .A(\parameter_B1_mul[7] ), .Y(n337) );
  INVX1 U7663 ( .A(\parameter_B2_mul[7] ), .Y(n328) );
  INVX1 U7664 ( .A(\parameter_A2_mul[7] ), .Y(n355) );
  INVX1 U7665 ( .A(\parameter_B0_mul[7] ), .Y(n346) );
  INVX1 U7666 ( .A(\parameter_A1_mul[7] ), .Y(n364) );
  INVX1 U7667 ( .A(\parameter_B1_mul[7] ), .Y(n338) );
  INVX1 U7668 ( .A(\parameter_B2_mul[7] ), .Y(n329) );
  INVX1 U7669 ( .A(\parameter_A1_mul[7] ), .Y(n365) );
  INVX1 U7670 ( .A(\parameter_A2_mul[7] ), .Y(n356) );
  INVX1 U7671 ( .A(\parameter_B0_mul[7] ), .Y(n347) );
endmodule

