
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_biquad_filter is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_biquad_filter;

library IEEE;

use IEEE.std_logic_1164.all;


use work.CONV_PACK_biquad_filter.all;

entity biquad_filter is

   port( clk, en, reset : in std_logic;  parameter_A1_mul, parameter_A1_div, 
         parameter_A2_mul, parameter_A2_div, parameter_B0_mul, parameter_B0_div
         , parameter_B1_mul, parameter_B1_div, parameter_B2_mul, 
         parameter_B2_div, input_signal : in std_logic_vector (7 downto 0);  
         output_signal : out std_logic_vector (7 downto 0);  change_input, 
         temporary_overflow : out std_logic);

end biquad_filter;

architecture SYN_flow_arch of biquad_filter is

   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A0, A1, B0, B1 : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR3XL
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI2BB1X1
      port( A0N, A1N, B0 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI2BB2X1
      port( B0, B1, A0N, A1N : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A0, A1, B0, B1 : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21XL
      port( A0, A1, B0 : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI221XL
      port( A0, A1, B0, B1, C0 : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2BX1
      port( AN, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI222XL
      port( A0, A1, B0, B1, C0, C1 : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI32X1
      port( A0, A1, A2, B0, B1 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2BX1
      port( AN, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3BX1
      port( AN, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2XL
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22XL
      port( A0, A1, B0, B1 : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2XL
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVXL
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFRXL
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRHQX1
      port( D, CK, RN : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSX1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2X4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal output_signal_7_port, output_signal_6_port, output_signal_5_port, 
      output_signal_4_port, output_signal_3_port, output_signal_2_port, 
      output_signal_1_port, n4673, input_previous_0_17_port, 
      input_previous_0_16_port, input_previous_0_15_port, 
      input_previous_0_14_port, input_previous_0_13_port, 
      input_previous_0_12_port, input_previous_0_11_port, 
      input_previous_0_10_port, input_previous_0_9_port, 
      input_previous_0_8_port, input_previous_0_7_port, input_previous_0_6_port
      , input_previous_0_5_port, input_previous_0_4_port, 
      input_previous_0_3_port, input_previous_0_2_port, input_previous_0_1_port
      , input_previous_1_17_port, input_previous_1_16_port, 
      input_previous_1_15_port, input_previous_1_14_port, 
      input_previous_1_13_port, input_previous_1_12_port, 
      input_previous_1_11_port, input_previous_1_10_port, 
      input_previous_1_9_port, input_previous_1_8_port, input_previous_1_7_port
      , input_previous_1_6_port, input_previous_1_5_port, 
      input_previous_1_4_port, input_previous_1_3_port, input_previous_1_2_port
      , input_previous_1_1_port, input_previous_2_17_port, 
      input_previous_2_16_port, input_previous_2_15_port, 
      input_previous_2_14_port, input_previous_2_13_port, 
      input_previous_2_12_port, input_previous_2_11_port, 
      input_previous_2_10_port, input_previous_2_9_port, 
      input_previous_2_8_port, input_previous_2_7_port, input_previous_2_6_port
      , input_previous_2_5_port, input_previous_2_4_port, 
      input_previous_2_3_port, input_previous_2_2_port, input_previous_2_1_port
      , output_previous_1_17_port, output_previous_1_16_port, 
      output_previous_1_15_port, output_previous_1_14_port, 
      output_previous_1_13_port, output_previous_1_12_port, 
      output_previous_1_11_port, output_previous_1_10_port, 
      output_previous_1_9_port, output_previous_1_8_port, 
      output_previous_2_17_port, output_previous_2_16_port, 
      output_previous_2_15_port, output_previous_2_14_port, 
      output_previous_2_13_port, output_previous_2_12_port, 
      output_previous_2_11_port, output_previous_2_10_port, 
      output_previous_2_9_port, output_previous_2_8_port, 
      output_previous_2_7_port, output_previous_2_6_port, 
      output_previous_2_5_port, output_previous_2_4_port, 
      output_previous_2_3_port, output_previous_2_2_port, 
      output_previous_2_1_port, results_b0_b1_17_port, results_b0_b1_16_port, 
      results_b0_b1_15_port, results_b0_b1_14_port, results_b0_b1_13_port, 
      results_b0_b1_12_port, results_b0_b1_11_port, results_b0_b1_10_port, 
      results_b0_b1_9_port, results_b0_b1_8_port, results_b0_b1_7_port, 
      results_b0_b1_6_port, results_b0_b1_5_port, results_b0_b1_4_port, 
      results_b0_b1_3_port, results_b0_b1_2_port, results_b0_b1_1_port, 
      results_b0_b1_0_port, results_b0_b1_b2_17_port, results_b0_b1_b2_16_port,
      results_b0_b1_b2_15_port, results_b0_b1_b2_14_port, 
      results_b0_b1_b2_13_port, results_b0_b1_b2_12_port, 
      results_b0_b1_b2_11_port, results_b0_b1_b2_10_port, 
      results_b0_b1_b2_9_port, results_b0_b1_b2_8_port, results_b0_b1_b2_7_port
      , results_b0_b1_b2_6_port, results_b0_b1_b2_5_port, 
      results_b0_b1_b2_4_port, results_b0_b1_b2_3_port, results_b0_b1_b2_2_port
      , results_b0_b1_b2_1_port, results_b0_b1_b2_0_port, results_a1_a2_17_port
      , results_a1_a2_16_port, results_a1_a2_15_port, results_a1_a2_14_port, 
      results_a1_a2_13_port, results_a1_a2_12_port, results_a1_a2_11_port, 
      results_a1_a2_10_port, results_a1_a2_9_port, results_a1_a2_8_port, 
      results_a1_a2_7_port, results_a1_a2_6_port, results_a1_a2_5_port, 
      results_a1_a2_4_port, results_a1_a2_3_port, results_a1_a2_2_port, 
      results_a1_a2_1_port, results_a1_a2_inv_17_port, 
      results_a1_a2_inv_16_port, results_a1_a2_inv_15_port, 
      results_a1_a2_inv_14_port, results_a1_a2_inv_13_port, 
      results_a1_a2_inv_12_port, results_a1_a2_inv_11_port, 
      results_a1_a2_inv_10_port, results_a1_a2_inv_9_port, 
      results_a1_a2_inv_8_port, results_a1_a2_inv_7_port, 
      results_a1_a2_inv_6_port, results_a1_a2_inv_5_port, 
      results_a1_a2_inv_4_port, results_a1_a2_inv_3_port, 
      results_a1_a2_inv_2_port, results_a1_a2_inv_1_port, 
      results_a1_a2_inv_0_port, output_contracterxn8, output_contracterxn7, 
      output_contracterxn6, output_contracterxn5, output_contracterxn4, 
      output_contracterxn3, output_contracterxn2, output_contracterxn1, 
      input_prev_0_registerxn20, input_prev_0_registerxn18, 
      input_prev_0_registerxn17, input_prev_0_registerxn16, 
      input_prev_0_registerxn15, input_prev_0_registerxn14, 
      input_prev_0_registerxn13, input_prev_0_registerxn12, 
      input_prev_0_registerxn11, input_prev_0_registerxn10, 
      input_prev_0_registerxn9, input_prev_0_registerxn8, 
      input_prev_0_registerxn7, input_prev_0_registerxn6, 
      input_prev_0_registerxn5, input_prev_0_registerxn4, 
      input_prev_0_registerxn3, input_prev_0_registerxn2, 
      input_times_b0_mul_componentxn108, input_times_b0_mul_componentxn107, 
      input_times_b0_mul_componentxn106, input_times_b0_mul_componentxn105, 
      input_times_b0_mul_componentxn104, input_times_b0_mul_componentxn103, 
      input_times_b0_mul_componentxn102, input_times_b0_mul_componentxn101, 
      input_times_b0_mul_componentxn100, input_times_b0_mul_componentxn99, 
      input_times_b0_mul_componentxn98, input_times_b0_mul_componentxn97, 
      input_times_b0_mul_componentxn96, input_times_b0_mul_componentxn95, 
      input_times_b0_mul_componentxn94, input_times_b0_mul_componentxn93, 
      input_times_b0_mul_componentxn92, input_times_b0_mul_componentxn91, 
      input_times_b0_mul_componentxn90, input_times_b0_mul_componentxn89, 
      input_times_b0_mul_componentxn88, input_times_b0_mul_componentxn87, 
      input_times_b0_mul_componentxn86, input_times_b0_mul_componentxn85, 
      input_times_b0_mul_componentxn84, input_times_b0_mul_componentxn83, 
      input_times_b0_mul_componentxn82, input_times_b0_mul_componentxn81, 
      input_times_b0_mul_componentxn80, input_times_b0_mul_componentxn79, 
      input_times_b0_mul_componentxn78, input_times_b0_mul_componentxn77, 
      input_times_b0_mul_componentxn76, input_times_b0_mul_componentxn75, 
      input_times_b0_mul_componentxn74, input_times_b0_mul_componentxn73, 
      input_times_b0_mul_componentxn72, input_times_b0_mul_componentxn71, 
      input_times_b0_mul_componentxn70, input_times_b0_mul_componentxn69, 
      input_times_b0_mul_componentxn68, input_times_b0_mul_componentxn67, 
      input_times_b0_mul_componentxn66, input_times_b0_mul_componentxn65, 
      input_times_b0_mul_componentxn64, input_times_b0_mul_componentxn63, 
      input_times_b0_mul_componentxn62, input_times_b0_mul_componentxn61, 
      input_times_b0_mul_componentxn60, input_times_b0_mul_componentxn59, 
      input_times_b0_mul_componentxn58, input_times_b0_mul_componentxn57, 
      input_times_b0_mul_componentxn56, 
      input_times_b0_mul_componentxunsigned_output_inverted_1_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_2_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_3_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_4_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_5_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_6_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_7_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_8_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_9_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_10_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_11_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_12_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_13_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_14_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_15_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_16_port, 
      input_times_b0_mul_componentxunsigned_output_inverted_17_port, 
      input_times_b0_mul_componentxunsigned_output_8, 
      input_times_b0_mul_componentxunsigned_output_9, 
      input_times_b0_mul_componentxunsigned_output_10, 
      input_times_b0_mul_componentxunsigned_output_11, 
      input_times_b0_mul_componentxunsigned_output_12, 
      input_times_b0_mul_componentxunsigned_output_13, 
      input_times_b0_mul_componentxunsigned_output_14, 
      input_times_b0_mul_componentxunsigned_output_15, 
      input_times_b0_mul_componentxunsigned_output_16, 
      input_times_b0_mul_componentxunsigned_output_17, 
      input_times_b0_mul_componentxinput_B_inverted_1_port, 
      input_times_b0_mul_componentxinput_B_inverted_2_port, 
      input_times_b0_mul_componentxinput_B_inverted_3_port, 
      input_times_b0_mul_componentxinput_B_inverted_4_port, 
      input_times_b0_mul_componentxinput_B_inverted_5_port, 
      input_times_b0_mul_componentxinput_B_inverted_6_port, 
      input_times_b0_mul_componentxinput_B_inverted_7_port, 
      input_times_b0_mul_componentxinput_B_inverted_8_port, 
      input_times_b0_mul_componentxinput_B_inverted_9_port, 
      input_times_b0_mul_componentxinput_B_inverted_10_port, 
      input_times_b0_mul_componentxinput_B_inverted_11_port, 
      input_times_b0_mul_componentxinput_B_inverted_12_port, 
      input_times_b0_mul_componentxinput_B_inverted_13_port, 
      input_times_b0_mul_componentxinput_B_inverted_14_port, 
      input_times_b0_mul_componentxinput_B_inverted_15_port, 
      input_times_b0_mul_componentxinput_B_inverted_16_port, 
      input_times_b0_mul_componentxinput_B_inverted_17_port, 
      input_times_b0_mul_componentxinput_A_inverted_0_port, 
      input_times_b0_mul_componentxinput_A_inverted_1_port, 
      input_times_b0_mul_componentxinput_A_inverted_2_port, 
      input_times_b0_mul_componentxinput_A_inverted_3_port, 
      input_times_b0_mul_componentxinput_A_inverted_4_port, 
      input_times_b0_mul_componentxinput_A_inverted_5_port, 
      input_times_b0_mul_componentxinput_A_inverted_6_port, 
      input_times_b0_mul_componentxinput_A_inverted_7_port, 
      input_times_b0_mul_componentxinput_A_inverted_8_port, 
      input_times_b0_mul_componentxinput_A_inverted_9_port, 
      input_times_b0_mul_componentxinput_A_inverted_10_port, 
      input_times_b0_mul_componentxinput_A_inverted_11_port, 
      input_times_b0_mul_componentxinput_A_inverted_12_port, 
      input_times_b0_mul_componentxinput_A_inverted_13_port, 
      input_times_b0_mul_componentxinput_A_inverted_14_port, 
      input_times_b0_mul_componentxinput_A_inverted_15_port, 
      input_times_b0_mul_componentxinput_A_inverted_16_port, 
      input_times_b0_mul_componentxinput_A_inverted_17_port, 
      input_times_b0_div_componentxn62, input_times_b0_div_componentxn61, 
      input_times_b0_div_componentxn60, input_times_b0_div_componentxn59, 
      input_times_b0_div_componentxn58, input_times_b0_div_componentxn57, 
      input_times_b0_div_componentxn56, input_times_b0_div_componentxn55, 
      input_times_b0_div_componentxn54, input_times_b0_div_componentxn53, 
      input_times_b0_div_componentxn52, input_times_b0_div_componentxn51, 
      input_times_b0_div_componentxn50, input_times_b0_div_componentxn49, 
      input_times_b0_div_componentxn48, input_times_b0_div_componentxn47, 
      input_times_b0_div_componentxn46, input_times_b0_div_componentxn45, 
      input_times_b0_div_componentxn44, input_times_b0_div_componentxn43, 
      input_times_b0_div_componentxn42, input_times_b0_div_componentxn41, 
      input_times_b0_div_componentxn40, input_times_b0_div_componentxn39, 
      input_times_b0_div_componentxn38, input_times_b0_div_componentxn37, 
      input_times_b0_div_componentxn36, input_times_b0_div_componentxn35, 
      input_times_b0_div_componentxn34, input_times_b0_div_componentxn33, 
      input_times_b0_div_componentxn32, input_times_b0_div_componentxn31, 
      input_times_b0_div_componentxn30, input_times_b0_div_componentxn29, 
      input_times_b0_div_componentxn28, input_times_b0_div_componentxn27, 
      input_times_b0_div_componentxn25, input_times_b0_div_componentxn24, 
      input_times_b0_div_componentxn21, input_times_b0_div_componentxn20, 
      input_times_b0_div_componentxn19, input_times_b0_div_componentxn18, 
      input_times_b0_div_componentxn17, input_times_b0_div_componentxn16, 
      input_times_b0_div_componentxn15, input_times_b0_div_componentxn14, 
      input_times_b0_div_componentxn13, input_times_b0_div_componentxn12, 
      input_times_b0_div_componentxn11, input_times_b0_div_componentxn10, 
      input_times_b0_div_componentxn9, input_times_b0_div_componentxn8, 
      input_times_b0_div_componentxn7, input_times_b0_div_componentxn6, 
      input_times_b0_div_componentxn5, input_times_b0_div_componentxn3, 
      input_times_b0_div_componentxoutput_sign_gated, 
      input_times_b0_div_componentxoutput_sign_gated_prev, 
      input_times_b0_div_componentxunsigned_B_17, 
      input_times_b0_div_componentxunsigned_A_17, 
      input_times_b0_div_componentxunsigned_output_inverted_0_port, 
      input_times_b0_div_componentxunsigned_output_inverted_1_port, 
      input_times_b0_div_componentxunsigned_output_inverted_2_port, 
      input_times_b0_div_componentxunsigned_output_inverted_3_port, 
      input_times_b0_div_componentxunsigned_output_inverted_4_port, 
      input_times_b0_div_componentxunsigned_output_inverted_5_port, 
      input_times_b0_div_componentxunsigned_output_inverted_6_port, 
      input_times_b0_div_componentxunsigned_output_inverted_7_port, 
      input_times_b0_div_componentxunsigned_output_inverted_8_port, 
      input_times_b0_div_componentxunsigned_output_inverted_9_port, 
      input_times_b0_div_componentxunsigned_output_inverted_10_port, 
      input_times_b0_div_componentxunsigned_output_inverted_11_port, 
      input_times_b0_div_componentxunsigned_output_inverted_12_port, 
      input_times_b0_div_componentxunsigned_output_inverted_13_port, 
      input_times_b0_div_componentxunsigned_output_inverted_14_port, 
      input_times_b0_div_componentxunsigned_output_inverted_15_port, 
      input_times_b0_div_componentxunsigned_output_inverted_16_port, 
      input_times_b0_div_componentxunsigned_output_inverted_17_port, 
      input_times_b0_div_componentxunsigned_output_1, 
      input_times_b0_div_componentxunsigned_output_2, 
      input_times_b0_div_componentxunsigned_output_3, 
      input_times_b0_div_componentxunsigned_output_4, 
      input_times_b0_div_componentxunsigned_output_5, 
      input_times_b0_div_componentxunsigned_output_6, 
      input_times_b0_div_componentxunsigned_output_7, 
      input_times_b0_div_componentxunsigned_output_8, 
      input_times_b0_div_componentxunsigned_output_9, 
      input_times_b0_div_componentxunsigned_output_10, 
      input_times_b0_div_componentxunsigned_output_11, 
      input_times_b0_div_componentxunsigned_output_12, 
      input_times_b0_div_componentxunsigned_output_13, 
      input_times_b0_div_componentxunsigned_output_14, 
      input_times_b0_div_componentxunsigned_output_15, 
      input_times_b0_div_componentxunsigned_output_16, 
      input_times_b0_div_componentxunsigned_output_17, 
      input_times_b0_div_componentxinput_B_inverted_1_port, 
      input_times_b0_div_componentxinput_B_inverted_2_port, 
      input_times_b0_div_componentxinput_B_inverted_3_port, 
      input_times_b0_div_componentxinput_B_inverted_4_port, 
      input_times_b0_div_componentxinput_B_inverted_5_port, 
      input_times_b0_div_componentxinput_B_inverted_6_port, 
      input_times_b0_div_componentxinput_B_inverted_7_port, 
      input_times_b0_div_componentxinput_B_inverted_8_port, 
      input_times_b0_div_componentxinput_B_inverted_9_port, 
      input_times_b0_div_componentxinput_B_inverted_10_port, 
      input_times_b0_div_componentxinput_B_inverted_11_port, 
      input_times_b0_div_componentxinput_B_inverted_12_port, 
      input_times_b0_div_componentxinput_B_inverted_13_port, 
      input_times_b0_div_componentxinput_B_inverted_14_port, 
      input_times_b0_div_componentxinput_B_inverted_15_port, 
      input_times_b0_div_componentxinput_B_inverted_16_port, 
      input_times_b0_div_componentxinput_B_inverted_17_port, 
      input_times_b0_div_componentxinput_A_inverted_1_port, 
      input_times_b0_div_componentxinput_A_inverted_2_port, 
      input_times_b0_div_componentxinput_A_inverted_3_port, 
      input_times_b0_div_componentxinput_A_inverted_4_port, 
      input_times_b0_div_componentxinput_A_inverted_5_port, 
      input_times_b0_div_componentxinput_A_inverted_6_port, 
      input_times_b0_div_componentxinput_A_inverted_7_port, 
      input_times_b0_div_componentxinput_A_inverted_8_port, 
      input_times_b0_div_componentxinput_A_inverted_9_port, 
      input_times_b0_div_componentxinput_A_inverted_10_port, 
      input_times_b0_div_componentxinput_A_inverted_11_port, 
      input_times_b0_div_componentxinput_A_inverted_12_port, 
      input_times_b0_div_componentxinput_A_inverted_13_port, 
      input_times_b0_div_componentxinput_A_inverted_14_port, 
      input_times_b0_div_componentxinput_A_inverted_15_port, 
      input_times_b0_div_componentxinput_A_inverted_16_port, 
      input_times_b0_div_componentxinput_A_inverted_17_port, 
      results_b0_b1_adderxn35, results_b0_b1_adderxn34, results_b0_b1_adderxn33
      , results_b0_b1_adderxn32, results_b0_b1_adderxn31, 
      results_b0_b1_adderxn30, results_b0_b1_adderxn29, results_b0_b1_adderxn28
      , results_b0_b1_adderxn27, results_b0_b1_adderxn26, 
      results_b0_b1_adderxn25, results_b0_b1_adderxn24, results_b0_b1_adderxn23
      , results_b0_b1_adderxn22, results_b0_b1_adderxn21, 
      results_b0_b1_adderxn20, results_b0_b1_adderxn19, results_b0_b1_adderxn17
      , results_b0_b1_adderxn16, results_b0_b1_adderxn15, 
      results_b0_b1_adderxn14, results_b0_b1_adderxn13, results_b0_b1_adderxn12
      , results_b0_b1_adderxn11, results_b0_b1_adderxn10, 
      results_b0_b1_adderxn9, results_b0_b1_adderxn8, results_b0_b1_adderxn7, 
      results_b0_b1_adderxn6, results_b0_b1_adderxn5, results_b0_b1_adderxn4, 
      results_b0_b1_adderxn3, results_b0_b1_adderxn2, 
      results_a1_a2_inv_inverterxn17, results_a1_a2_inv_inverterxn15, 
      results_a1_a2_inv_inverterxn13, results_a1_a2_inv_inverterxn12, 
      results_a1_a2_inv_inverterxn11, results_a1_a2_inv_inverterxn10, 
      results_a1_a2_inv_inverterxn9, results_a1_a2_inv_inverterxn8, 
      results_a1_a2_inv_inverterxn6, results_a1_a2_inv_inverterxn4, 
      results_a1_a2_inv_inverterxn2, clock_chopper_and_divisionxn49, 
      clock_chopper_and_divisionxn47, clock_chopper_and_divisionxn46, 
      clock_chopper_and_divisionxn45, clock_chopper_and_divisionxn44, 
      clock_chopper_and_divisionxn43, clock_chopper_and_divisionxn42, 
      clock_chopper_and_divisionxn41, clock_chopper_and_divisionxn40, 
      clock_chopper_and_divisionxn39, clock_chopper_and_divisionxn38, 
      clock_chopper_and_divisionxn37, clock_chopper_and_divisionxn36, 
      clock_chopper_and_divisionxn35, clock_chopper_and_divisionxn34, 
      clock_chopper_and_divisionxn33, clock_chopper_and_divisionxn32, 
      clock_chopper_and_divisionxn31, clock_chopper_and_divisionxn30, 
      clock_chopper_and_divisionxn29, clock_chopper_and_divisionxn28, 
      clock_chopper_and_divisionxn27, clock_chopper_and_divisionxn26, 
      clock_chopper_and_divisionxdivision_ring_0_port, 
      clock_chopper_and_divisionxdivision_ring_1_port, 
      clock_chopper_and_divisionxdivision_ring_2_port, 
      clock_chopper_and_divisionxdivision_ring_3_port, 
      clock_chopper_and_divisionxdivision_ring_4_port, 
      clock_chopper_and_divisionxdivision_ring_5_port, 
      clock_chopper_and_divisionxdivision_ring_6_port, 
      clock_chopper_and_divisionxdivision_ring_7_port, 
      clock_chopper_and_divisionxdivision_ring_8_port, 
      clock_chopper_and_divisionxdivision_ring_9_port, 
      clock_chopper_and_divisionxdivision_ring_10_port, 
      clock_chopper_and_divisionxdivision_ring_11_port, 
      clock_chopper_and_divisionxdivision_ring_12_port, 
      clock_chopper_and_divisionxdivision_ring_13_port, 
      clock_chopper_and_divisionxdivision_ring_14_port, 
      clock_chopper_and_divisionxdivision_ring_15_port, 
      clock_chopper_and_divisionxdivision_ring_16_port, 
      clock_chopper_and_divisionxdivision_ring_17_port, 
      clock_chopper_and_divisionxdivision_ring_18_port, 
      clock_chopper_and_divisionxdivision_ring_19_port, 
      clock_chopper_and_divisionxdivision_ring_20_port, 
      clock_chopper_and_divisionxdivision_ring_21_port, 
      input_times_b0_mul_componentxUMxsecond_vector_7_port, 
      input_times_b0_mul_componentxUMxsecond_vector_8_port, 
      input_times_b0_mul_componentxUMxsecond_vector_9_port, 
      input_times_b0_mul_componentxUMxsecond_vector_10_port, 
      input_times_b0_mul_componentxUMxsecond_vector_11_port, 
      input_times_b0_mul_componentxUMxsecond_vector_12_port, 
      input_times_b0_mul_componentxUMxsecond_vector_13_port, 
      input_times_b0_mul_componentxUMxsecond_vector_14_port, 
      input_times_b0_mul_componentxUMxsecond_vector_15_port, 
      input_times_b0_mul_componentxUMxsecond_vector_16_port, 
      input_times_b0_mul_componentxUMxsecond_vector_17_port, 
      input_times_b0_mul_componentxUMxfirst_vector_0_port, 
      input_times_b0_mul_componentxUMxfirst_vector_1_port, 
      input_times_b0_mul_componentxUMxfirst_vector_2_port, 
      input_times_b0_mul_componentxUMxfirst_vector_3_port, 
      input_times_b0_mul_componentxUMxfirst_vector_4_port, 
      input_times_b0_mul_componentxUMxfirst_vector_5_port, 
      input_times_b0_mul_componentxUMxfirst_vector_6_port, 
      input_times_b0_mul_componentxUMxfirst_vector_7_port, 
      input_times_b0_mul_componentxUMxfirst_vector_8_port, 
      input_times_b0_mul_componentxUMxfirst_vector_9_port, 
      input_times_b0_mul_componentxUMxfirst_vector_10_port, 
      input_times_b0_mul_componentxUMxfirst_vector_11_port, 
      input_times_b0_mul_componentxUMxfirst_vector_12_port, 
      input_times_b0_mul_componentxUMxfirst_vector_13_port, 
      input_times_b0_mul_componentxUMxfirst_vector_14_port, 
      input_times_b0_mul_componentxUMxfirst_vector_15_port, 
      input_times_b0_mul_componentxUMxsum_layer5_128315744_128315968_128316136,
      input_times_b0_mul_componentxUMxsum_layer5_128315464_128315632_128315800,
      input_times_b0_mul_componentxUMxsum_layer5_128220800_128221024_128221136,
      input_times_b0_mul_componentxUMxsum_layer5_128220688_128220856_128220968,
      input_times_b0_mul_componentxUMxsum_layer5_128126256_128220520_128220744,
      input_times_b0_mul_componentxUMxsum_layer5_128125920_128220352_128220576,
      input_times_b0_mul_componentxUMxsum_layer5_128125584_128220184_128220408,
      input_times_b0_mul_componentxUMxsum_layer5_128125248_128219960_128220240,
      input_times_b0_mul_componentxUMxcarry_layer5_128219792_128220016, 
      input_times_b0_mul_componentxUMxsum_layer5_128219792_128220016, 
      input_times_b0_mul_componentxUMxcarry_layer5_128219624_128219848, 
      input_times_b0_mul_componentxUMxsum_layer5_128219624_128219848, 
      input_times_b0_mul_componentxUMxcarry_layer5_128219456_128219680, 
      input_times_b0_mul_componentxUMxsum_layer5_128219456_128219680, 
      input_times_b0_mul_componentxUMxcarry_layer5_128219288_128219512, 
      input_times_b0_mul_componentxUMxsum_layer5_128219288_128219512, 
      input_times_b0_mul_componentxUMxcarry_layer5_128219120_128219344, 
      input_times_b0_mul_componentxUMxsum_layer4_128238312_128238424_128238592,
      input_times_b0_mul_componentxUMxsum_layer4_128237752_128237976_128238144,
      input_times_b0_mul_componentxUMxsum_layer4_128237920_128238088, 
      input_times_b0_mul_componentxUMxsum_layer4_128126760_128237640_128237808,
      input_times_b0_mul_componentxUMxcarry_layer4_128126816_128126928, 
      input_times_b0_mul_componentxUMxsum_layer4_128126816_128126928, 
      input_times_b0_mul_componentxUMxsum_layer4_128263168_128126424_128126648,
      input_times_b0_mul_componentxUMxcarry_layer4_128126480_128126592, 
      input_times_b0_mul_componentxUMxsum_layer4_128126480_128126592, 
      input_times_b0_mul_componentxUMxsum_layer4_128262496_128126088_128126312,
      input_times_b0_mul_componentxUMxsum_layer4_128125752_128125976_128126144,
      input_times_b0_mul_componentxUMxsum_layer4_128125416_128125640_128125808,
      input_times_b0_mul_componentxUMxsum_layer4_128125080_128125304_128125472,
      input_times_b0_mul_componentxUMxsum_layer4_128124744_128124968_128125136,
      input_times_b0_mul_componentxUMxsum_layer4_128124632_128124800_128124912,
      input_times_b0_mul_componentxUMxsum_layer4_128247456_128124464_128124688,
      input_times_b0_mul_componentxUMxsum_layer4_128247120_128124240_128124520,
      input_times_b0_mul_componentxUMxcarry_layer4_128124072_128124296, 
      input_times_b0_mul_componentxUMxsum_layer4_128124072_128124296, 
      input_times_b0_mul_componentxUMxcarry_layer4_128123904_128124128, 
      input_times_b0_mul_componentxUMxsum_layer4_128123904_128124128, 
      input_times_b0_mul_componentxUMxcarry_layer4_128123792_128123960, 
      input_times_b0_mul_componentxUMxsum_layer3_128264344_128264512, 
      input_times_b0_mul_componentxUMxsum_layer3_128263896_128264064_128264176,
      input_times_b0_mul_componentxUMxsum_layer3_128263336_128263560_128263728,
      input_times_b0_mul_componentxUMxcarry_layer3_128263672_128263840, 
      input_times_b0_mul_componentxUMxsum_layer3_128263672_128263840, 
      input_times_b0_mul_componentxUMxsum_layer3_128263224_128263392_128263504,
      input_times_b0_mul_componentxUMxsum_layer3_128262664_128262888_128263056,
      input_times_b0_mul_componentxUMxsum_layer3_128262720_128262832_128263000,
      input_times_b0_mul_componentxUMxsum_layer3_128262216_128262384_128262552,
      input_times_b0_mul_componentxUMxsum_layer3_128249696_128249808_128262328,
      input_times_b0_mul_componentxUMxsum_layer3_128197128_128249304_128249528,
      input_times_b0_mul_componentxUMxsum_layer3_128249360_128249472_128249640,
      input_times_b0_mul_componentxUMxsum_layer3_128248800_128249024_128249192,
      input_times_b0_mul_componentxUMxsum_layer3_128248856_128248968_128249136,
      input_times_b0_mul_componentxUMxsum_layer3_128248296_128248520_128248688,
      input_times_b0_mul_componentxUMxcarry_layer3_128248464_128248632, 
      input_times_b0_mul_componentxUMxsum_layer3_128248464_128248632, 
      input_times_b0_mul_componentxUMxsum_layer3_128247960_128248184_128248352,
      input_times_b0_mul_componentxUMxcarry_layer3_128248016_128248128, 
      input_times_b0_mul_componentxUMxsum_layer3_128248016_128248128, 
      input_times_b0_mul_componentxUMxsum_layer3_128222880_128247624_128247848,
      input_times_b0_mul_componentxUMxcarry_layer3_128247680_128247792, 
      input_times_b0_mul_componentxUMxsum_layer3_128247680_128247792, 
      input_times_b0_mul_componentxUMxsum_layer3_128222208_128247288_128247512,
      input_times_b0_mul_componentxUMxsum_layer3_128246952_128247176_128247344,
      input_times_b0_mul_componentxUMxsum_layer3_128246616_128246840_128247008,
      input_times_b0_mul_componentxUMxsum_layer3_128246504_128246672_128246784,
      input_times_b0_mul_componentxUMxsum_layer3_127827080_128246280_128246560,
      input_times_b0_mul_componentxUMxcarry_layer3_128246112_128246336, 
      input_times_b0_mul_componentxUMxsum_layer3_128246112_128246336, 
      input_times_b0_mul_componentxUMxcarry_layer3_128246000_128246168, 
      input_times_b0_mul_componentxUMxsum_layer2_128199816_128200040_128199984,
      input_times_b0_mul_componentxUMxsum_layer2_128199368_128199480_128199648,
      input_times_b0_mul_componentxUMxsum_layer2_128198864_128199032_128199200,
      input_times_b0_mul_componentxUMxsum_layer2_128198304_128198528_128198696,
      input_times_b0_mul_componentxUMxcarry_layer2_128198976_128199144, 
      input_times_b0_mul_componentxUMxsum_layer2_128198976_128199144, 
      input_times_b0_mul_componentxUMxsum_layer2_128198472_128198640_128198808,
      input_times_b0_mul_componentxUMxsum_layer2_128198080_128198192_128198360,
      input_times_b0_mul_componentxUMxsum_layer2_128197464_128197688_128197856,
      input_times_b0_mul_componentxUMxcarry_layer2_128198024_128197968, 
      input_times_b0_mul_componentxUMxsum_layer2_128198024_128197968, 
      input_times_b0_mul_componentxUMxsum_layer2_128197520_128197632_128197800,
      input_times_b0_mul_componentxUMxsum_layer2_128197016_128197240_128197352,
      input_times_b0_mul_componentxUMxsum_layer2_127627392_128196680_128196848,
      input_times_b0_mul_componentxUMxa15_and_b0, 
      input_times_b0_mul_componentxUMxsum_layer2_128196792_128196960_128197184,
      input_times_b0_mul_componentxUMxsum_layer2_128224952_128225120_128225232,
      input_times_b0_mul_componentxUMxsum_layer2_128224392_128224616_128224784,
      input_times_b0_mul_componentxUMxsum_layer2_128224728_128224896_128225064,
      input_times_b0_mul_componentxUMxsum_layer2_128224280_128224448_128224560,
      input_times_b0_mul_componentxUMxsum_layer2_128223720_128223944_128224168,
      input_times_b0_mul_componentxUMxsum_layer2_128223888_128224112_128224056,
      input_times_b0_mul_componentxUMxsum_layer2_128223440_128223608_128223776,
      input_times_b0_mul_componentxUMxsum_layer2_127715424_128223048_128223272,
      input_times_b0_mul_componentxUMxa12_and_b0, 
      input_times_b0_mul_componentxUMxcarry_layer2_128223384_128223552, 
      input_times_b0_mul_componentxUMxsum_layer2_128223384_128223552, 
      input_times_b0_mul_componentxUMxsum_layer2_128222936_128223104_128223216,
      input_times_b0_mul_componentxUMxsum_layer2_128222376_128222600_128222768,
      input_times_b0_mul_componentxUMxsum_layer2_128222432_128222544_128222712,
      input_times_b0_mul_componentxUMxsum_layer2_128221872_128222096_128222264,
      input_times_b0_mul_componentxUMxsum_layer2_128221760_128221928_128222040,
      input_times_b0_mul_componentxUMxsum_layer2_127635584_128221368_128221592,
      input_times_b0_mul_componentxUMxa9_and_b0, 
      input_times_b0_mul_componentxUMxsum_layer2_128221424_128221536_128221704,
      input_times_b0_mul_componentxUMxsum_layer2_127827584_127827808_128221256,
      input_times_b0_mul_componentxUMxcarry_layer2_127827752_127827920, 
      input_times_b0_mul_componentxUMxsum_layer2_127827752_127827920, 
      input_times_b0_mul_componentxUMxsum_layer2_127827248_127827472_127827640,
      input_times_b0_mul_componentxUMxcarry_layer2_127827304_127827416, 
      input_times_b0_mul_componentxUMxsum_layer2_127827304_127827416, 
      input_times_b0_mul_componentxUMxsum_layer2_127731808_127826912_127827136,
      input_times_b0_mul_componentxUMxa6_and_b0, 
      input_times_b0_mul_componentxUMxsum_layer2_127826576_127826800_127826968,
      input_times_b0_mul_componentxUMxsum_layer2_127826464_127826632_127826744,
      input_times_b0_mul_componentxUMxsum_layer2_127672448_127826240_127826520,
      input_times_b0_mul_componentxUMxa3_and_b0, 
      input_times_b0_mul_componentxUMxcarry_layer2_127826128_127826296, 
      input_times_b0_mul_componentxUMxsum_layer1_127627616_127629520_127824000,
      input_times_b0_mul_componentxUMxa17_and_b0, 
      input_times_b0_mul_componentxUMxa16_and_b1, 
      input_times_b0_mul_componentxUMxa15_and_b2, 
      input_times_b0_mul_componentxUMxsum_layer1_127715984_127849024_127850928,
      input_times_b0_mul_componentxUMxa14_and_b3, 
      input_times_b0_mul_componentxUMxa13_and_b4, 
      input_times_b0_mul_componentxUMxa12_and_b5, 
      input_times_b0_mul_componentxUMxsum_layer1_127636480_127638384_127714080,
      input_times_b0_mul_componentxUMxa11_and_b6, 
      input_times_b0_mul_componentxUMxa10_and_b7, 
      input_times_b0_mul_componentxUMxa9_and_b8, 
      input_times_b0_mul_componentxUMxsum_layer1_127733040_127722720_127724624,
      input_times_b0_mul_componentxUMxa8_and_b9, 
      input_times_b0_mul_componentxUMxa7_and_b10, 
      input_times_b0_mul_componentxUMxa6_and_b11, 
      input_times_b0_mul_componentxUMxsum_layer1_127674016_127675920_127731136,
      input_times_b0_mul_componentxUMxa5_and_b12, 
      input_times_b0_mul_componentxUMxa4_and_b13, 
      input_times_b0_mul_componentxUMxa3_and_b14, 
      input_times_b0_mul_componentxUMxsum_layer1_127832016_127846272_127848176,
      input_times_b0_mul_componentxUMxa2_and_b15, 
      input_times_b0_mul_componentxUMxa1_and_b16, 
      input_times_b0_mul_componentxUMxa0_and_b17, 
      input_times_b0_mul_componentxUMxcarry_layer1_127627504_127629408, 
      input_times_b0_mul_componentxUMxsum_layer1_127627504_127629408, 
      input_times_b0_mul_componentxUMxa16_and_b0, 
      input_times_b0_mul_componentxUMxa15_and_b1, 
      input_times_b0_mul_componentxUMxsum_layer1_127715872_127848912_127850816,
      input_times_b0_mul_componentxUMxa14_and_b2, 
      input_times_b0_mul_componentxUMxa13_and_b3, 
      input_times_b0_mul_componentxUMxa12_and_b4, 
      input_times_b0_mul_componentxUMxsum_layer1_127636368_127638272_127713968,
      input_times_b0_mul_componentxUMxa11_and_b5, 
      input_times_b0_mul_componentxUMxa10_and_b6, 
      input_times_b0_mul_componentxUMxa9_and_b7, 
      input_times_b0_mul_componentxUMxsum_layer1_127732928_127722608_127724512,
      input_times_b0_mul_componentxUMxa8_and_b8, 
      input_times_b0_mul_componentxUMxa7_and_b9, 
      input_times_b0_mul_componentxUMxa6_and_b10, 
      input_times_b0_mul_componentxUMxsum_layer1_127673904_127675808_127731024,
      input_times_b0_mul_componentxUMxa5_and_b11, 
      input_times_b0_mul_componentxUMxa4_and_b12, 
      input_times_b0_mul_componentxUMxa3_and_b13, 
      input_times_b0_mul_componentxUMxsum_layer1_127831904_127846160_127848064,
      input_times_b0_mul_componentxUMxa2_and_b14, 
      input_times_b0_mul_componentxUMxa1_and_b15, 
      input_times_b0_mul_componentxUMxa0_and_b16, 
      input_times_b0_mul_componentxUMxsum_layer1_127715760_127848800_127850704,
      input_times_b0_mul_componentxUMxa14_and_b1, 
      input_times_b0_mul_componentxUMxa13_and_b2, 
      input_times_b0_mul_componentxUMxa12_and_b3, 
      input_times_b0_mul_componentxUMxsum_layer1_127636256_127638160_127713856,
      input_times_b0_mul_componentxUMxa11_and_b4, 
      input_times_b0_mul_componentxUMxa10_and_b5, 
      input_times_b0_mul_componentxUMxa9_and_b6, 
      input_times_b0_mul_componentxUMxsum_layer1_127732816_127722496_127724400,
      input_times_b0_mul_componentxUMxa8_and_b7, 
      input_times_b0_mul_componentxUMxa7_and_b8, 
      input_times_b0_mul_componentxUMxa6_and_b9, 
      input_times_b0_mul_componentxUMxsum_layer1_127673792_127675696_127730912,
      input_times_b0_mul_componentxUMxa5_and_b10, 
      input_times_b0_mul_componentxUMxa4_and_b11, 
      input_times_b0_mul_componentxUMxa3_and_b12, 
      input_times_b0_mul_componentxUMxsum_layer1_127831792_127846048_127847952,
      input_times_b0_mul_componentxUMxa2_and_b13, 
      input_times_b0_mul_componentxUMxa1_and_b14, 
      input_times_b0_mul_componentxUMxa0_and_b15, 
      input_times_b0_mul_componentxUMxsum_layer1_127715648_127848688_127850592,
      input_times_b0_mul_componentxUMxa14_and_b0, 
      input_times_b0_mul_componentxUMxa13_and_b1, 
      input_times_b0_mul_componentxUMxa12_and_b2, 
      input_times_b0_mul_componentxUMxsum_layer1_127636144_127638048_127713744,
      input_times_b0_mul_componentxUMxa11_and_b3, 
      input_times_b0_mul_componentxUMxa10_and_b4, 
      input_times_b0_mul_componentxUMxa9_and_b5, 
      input_times_b0_mul_componentxUMxsum_layer1_127732704_127722384_127724288,
      input_times_b0_mul_componentxUMxa8_and_b6, 
      input_times_b0_mul_componentxUMxa7_and_b7, 
      input_times_b0_mul_componentxUMxa6_and_b8, 
      input_times_b0_mul_componentxUMxsum_layer1_127673680_127675584_127730800,
      input_times_b0_mul_componentxUMxa5_and_b9, 
      input_times_b0_mul_componentxUMxa4_and_b10, 
      input_times_b0_mul_componentxUMxa3_and_b11, 
      input_times_b0_mul_componentxUMxsum_layer1_127831680_127845936_127847840,
      input_times_b0_mul_componentxUMxa2_and_b12, 
      input_times_b0_mul_componentxUMxa1_and_b13, 
      input_times_b0_mul_componentxUMxa0_and_b14, 
      input_times_b0_mul_componentxUMxcarry_layer1_127715536_127848576, 
      input_times_b0_mul_componentxUMxsum_layer1_127715536_127848576, 
      input_times_b0_mul_componentxUMxa13_and_b0, 
      input_times_b0_mul_componentxUMxa12_and_b1, 
      input_times_b0_mul_componentxUMxsum_layer1_127636032_127637936_127713632,
      input_times_b0_mul_componentxUMxa11_and_b2, 
      input_times_b0_mul_componentxUMxa10_and_b3, 
      input_times_b0_mul_componentxUMxa9_and_b4, 
      input_times_b0_mul_componentxUMxsum_layer1_127732592_127722272_127724176,
      input_times_b0_mul_componentxUMxa8_and_b5, 
      input_times_b0_mul_componentxUMxa7_and_b6, 
      input_times_b0_mul_componentxUMxa6_and_b7, 
      input_times_b0_mul_componentxUMxsum_layer1_127673568_127675472_127730688,
      input_times_b0_mul_componentxUMxa5_and_b8, 
      input_times_b0_mul_componentxUMxa4_and_b9, 
      input_times_b0_mul_componentxUMxa3_and_b10, 
      input_times_b0_mul_componentxUMxsum_layer1_127831568_127845824_127847728,
      input_times_b0_mul_componentxUMxa2_and_b11, 
      input_times_b0_mul_componentxUMxa1_and_b12, 
      input_times_b0_mul_componentxUMxa0_and_b13, 
      input_times_b0_mul_componentxUMxsum_layer1_127635920_127637824_127713520,
      input_times_b0_mul_componentxUMxa11_and_b1, 
      input_times_b0_mul_componentxUMxa10_and_b2, 
      input_times_b0_mul_componentxUMxa9_and_b3, 
      input_times_b0_mul_componentxUMxsum_layer1_127732480_127722160_127724064,
      input_times_b0_mul_componentxUMxa8_and_b4, 
      input_times_b0_mul_componentxUMxa7_and_b5, 
      input_times_b0_mul_componentxUMxa6_and_b6, 
      input_times_b0_mul_componentxUMxsum_layer1_127673456_127675360_127730576,
      input_times_b0_mul_componentxUMxa5_and_b7, 
      input_times_b0_mul_componentxUMxa4_and_b8, 
      input_times_b0_mul_componentxUMxa3_and_b9, 
      input_times_b0_mul_componentxUMxsum_layer1_127831456_127845712_127847616,
      input_times_b0_mul_componentxUMxa2_and_b10, 
      input_times_b0_mul_componentxUMxa1_and_b11, 
      input_times_b0_mul_componentxUMxa0_and_b12, 
      input_times_b0_mul_componentxUMxsum_layer1_127635808_127637712_127713408,
      input_times_b0_mul_componentxUMxa11_and_b0, 
      input_times_b0_mul_componentxUMxa10_and_b1, 
      input_times_b0_mul_componentxUMxa9_and_b2, 
      input_times_b0_mul_componentxUMxsum_layer1_127732368_127722048_127723952,
      input_times_b0_mul_componentxUMxa8_and_b3, 
      input_times_b0_mul_componentxUMxa7_and_b4, 
      input_times_b0_mul_componentxUMxa6_and_b5, 
      input_times_b0_mul_componentxUMxsum_layer1_127673344_127675248_127730464,
      input_times_b0_mul_componentxUMxa5_and_b6, 
      input_times_b0_mul_componentxUMxa4_and_b7, 
      input_times_b0_mul_componentxUMxa3_and_b8, 
      input_times_b0_mul_componentxUMxsum_layer1_127831344_127845600_127847504,
      input_times_b0_mul_componentxUMxa2_and_b9, 
      input_times_b0_mul_componentxUMxa1_and_b10, 
      input_times_b0_mul_componentxUMxa0_and_b11, 
      input_times_b0_mul_componentxUMxcarry_layer1_127635696_127637600, 
      input_times_b0_mul_componentxUMxsum_layer1_127635696_127637600, 
      input_times_b0_mul_componentxUMxa10_and_b0, 
      input_times_b0_mul_componentxUMxa9_and_b1, 
      input_times_b0_mul_componentxUMxsum_layer1_127732256_127721936_127723840,
      input_times_b0_mul_componentxUMxa8_and_b2, 
      input_times_b0_mul_componentxUMxa7_and_b3, 
      input_times_b0_mul_componentxUMxa6_and_b4, 
      input_times_b0_mul_componentxUMxsum_layer1_127673232_127675136_127730352,
      input_times_b0_mul_componentxUMxa5_and_b5, 
      input_times_b0_mul_componentxUMxa4_and_b6, 
      input_times_b0_mul_componentxUMxa3_and_b7, 
      input_times_b0_mul_componentxUMxsum_layer1_127831232_127845488_127847392,
      input_times_b0_mul_componentxUMxa2_and_b8, 
      input_times_b0_mul_componentxUMxa1_and_b9, 
      input_times_b0_mul_componentxUMxa0_and_b10, 
      input_times_b0_mul_componentxUMxsum_layer1_127732144_127721824_127723728,
      input_times_b0_mul_componentxUMxa8_and_b1, 
      input_times_b0_mul_componentxUMxa7_and_b2, 
      input_times_b0_mul_componentxUMxa6_and_b3, 
      input_times_b0_mul_componentxUMxsum_layer1_127673120_127675024_127730240,
      input_times_b0_mul_componentxUMxa5_and_b4, 
      input_times_b0_mul_componentxUMxa4_and_b5, 
      input_times_b0_mul_componentxUMxa3_and_b6, 
      input_times_b0_mul_componentxUMxsum_layer1_127831120_127845376_127847280,
      input_times_b0_mul_componentxUMxa2_and_b7, 
      input_times_b0_mul_componentxUMxa1_and_b8, 
      input_times_b0_mul_componentxUMxa0_and_b9, 
      input_times_b0_mul_componentxUMxsum_layer1_127732032_127721712_127723616,
      input_times_b0_mul_componentxUMxa8_and_b0, 
      input_times_b0_mul_componentxUMxa7_and_b1, 
      input_times_b0_mul_componentxUMxa6_and_b2, 
      input_times_b0_mul_componentxUMxsum_layer1_127673008_127674912_127730128,
      input_times_b0_mul_componentxUMxa5_and_b3, 
      input_times_b0_mul_componentxUMxa4_and_b4, 
      input_times_b0_mul_componentxUMxa3_and_b5, 
      input_times_b0_mul_componentxUMxsum_layer1_127831008_127845264_127847168,
      input_times_b0_mul_componentxUMxa2_and_b6, 
      input_times_b0_mul_componentxUMxa1_and_b7, 
      input_times_b0_mul_componentxUMxa0_and_b8, 
      input_times_b0_mul_componentxUMxcarry_layer1_127731920_127721600, 
      input_times_b0_mul_componentxUMxsum_layer1_127731920_127721600, 
      input_times_b0_mul_componentxUMxa7_and_b0, 
      input_times_b0_mul_componentxUMxa6_and_b1, 
      input_times_b0_mul_componentxUMxsum_layer1_127672896_127674800_127730016,
      input_times_b0_mul_componentxUMxa5_and_b2, 
      input_times_b0_mul_componentxUMxa4_and_b3, 
      input_times_b0_mul_componentxUMxa3_and_b4, 
      input_times_b0_mul_componentxUMxsum_layer1_127830896_127845152_127847056,
      input_times_b0_mul_componentxUMxa2_and_b5, 
      input_times_b0_mul_componentxUMxa1_and_b6, 
      input_times_b0_mul_componentxUMxa0_and_b7, 
      input_times_b0_mul_componentxUMxsum_layer1_127672784_127674688_127729904,
      input_times_b0_mul_componentxUMxa5_and_b1, 
      input_times_b0_mul_componentxUMxa4_and_b2, 
      input_times_b0_mul_componentxUMxa3_and_b3, 
      input_times_b0_mul_componentxUMxsum_layer1_127830784_127845040_127846944,
      input_times_b0_mul_componentxUMxa2_and_b4, 
      input_times_b0_mul_componentxUMxa1_and_b5, 
      input_times_b0_mul_componentxUMxa0_and_b6, 
      input_times_b0_mul_componentxUMxsum_layer1_127672672_127674576_127729792,
      input_times_b0_mul_componentxUMxa5_and_b0, 
      input_times_b0_mul_componentxUMxa4_and_b1, 
      input_times_b0_mul_componentxUMxa3_and_b2, 
      input_times_b0_mul_componentxUMxsum_layer1_127830672_127844928_127846832,
      input_times_b0_mul_componentxUMxa2_and_b3, 
      input_times_b0_mul_componentxUMxa1_and_b4, 
      input_times_b0_mul_componentxUMxa0_and_b5, 
      input_times_b0_mul_componentxUMxcarry_layer1_127672560_127674464, 
      input_times_b0_mul_componentxUMxsum_layer1_127672560_127674464, 
      input_times_b0_mul_componentxUMxa4_and_b0, 
      input_times_b0_mul_componentxUMxa3_and_b1, 
      input_times_b0_mul_componentxUMxsum_layer1_127830560_127844816_127846720,
      input_times_b0_mul_componentxUMxa2_and_b2, 
      input_times_b0_mul_componentxUMxa1_and_b3, 
      input_times_b0_mul_componentxUMxa0_and_b4, 
      input_times_b0_mul_componentxUMxsum_layer1_127830448_127844704_127846608,
      input_times_b0_mul_componentxUMxa2_and_b1, 
      input_times_b0_mul_componentxUMxa1_and_b2, 
      input_times_b0_mul_componentxUMxa0_and_b3, 
      input_times_b0_mul_componentxUMxsum_layer1_127830336_127844592_127846496,
      input_times_b0_mul_componentxUMxa2_and_b0, 
      input_times_b0_mul_componentxUMxa1_and_b1, 
      input_times_b0_mul_componentxUMxa0_and_b2, 
      input_times_b0_mul_componentxUMxcarry_layer1_127830168_127844480, 
      input_times_b0_mul_componentxUMxa1_and_b0, 
      input_times_b0_mul_componentxUMxa0_and_b1, 
      input_times_b0_div_componentxUDxn19, input_times_b0_div_componentxUDxn18,
      input_times_b0_div_componentxUDxn17, input_times_b0_div_componentxUDxn16,
      input_times_b0_div_componentxUDxn15, input_times_b0_div_componentxUDxn14,
      input_times_b0_div_componentxUDxn13, input_times_b0_div_componentxUDxn12,
      input_times_b0_div_componentxUDxn11, input_times_b0_div_componentxUDxn10,
      input_times_b0_div_componentxUDxn9, input_times_b0_div_componentxUDxn8, 
      input_times_b0_div_componentxUDxn7, input_times_b0_div_componentxUDxn6, 
      input_times_b0_div_componentxUDxn5, input_times_b0_div_componentxUDxn4, 
      input_times_b0_div_componentxUDxn3, input_times_b0_div_componentxUDxn1, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_0_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_1_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_2_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_3_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_4_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_5_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_6_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_7_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_8_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_9_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_10_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_11_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_12_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_13_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_14_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_15_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_16_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_17_port, 
      input_times_b0_div_componentxUDxreadiness_propagation_vector_18_port, 
      input_times_b0_div_componentxUDxis_less_than, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_0_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_1_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_2_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_3_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_4_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_5_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_6_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_7_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_8_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_9_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_10_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_11_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_12_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_13_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_14_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_15_port, 
      input_times_b0_div_componentxUDxsubstraction_result_too_long_16_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_1_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_2_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_3_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_4_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_5_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_6_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_7_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_8_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_9_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_10_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_11_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_12_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_13_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_14_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_15_port, 
      input_times_b0_div_componentxUDxsub_ready_negative_divisor_16_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_0_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_1_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_2_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_3_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_4_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_5_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_6_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_7_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_8_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_9_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_10_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_11_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_12_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_13_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_14_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_15_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_16_port, 
      input_times_b0_div_componentxUDxquotient_not_gated_17_port, 
      input_times_b0_div_componentxUDxcentral_parallel_output_0, 
      input_times_b0_div_componentxUDxcentral_parallel_output_1, 
      input_times_b0_div_componentxUDxcentral_parallel_output_2, 
      input_times_b0_div_componentxUDxcentral_parallel_output_3, 
      input_times_b0_div_componentxUDxcentral_parallel_output_4, 
      input_times_b0_div_componentxUDxcentral_parallel_output_5, 
      input_times_b0_div_componentxUDxcentral_parallel_output_6, 
      input_times_b0_div_componentxUDxcentral_parallel_output_7, 
      input_times_b0_div_componentxUDxcentral_parallel_output_8, 
      input_times_b0_div_componentxUDxcentral_parallel_output_9, 
      input_times_b0_div_componentxUDxcentral_parallel_output_10, 
      input_times_b0_div_componentxUDxcentral_parallel_output_11, 
      input_times_b0_div_componentxUDxcentral_parallel_output_12, 
      input_times_b0_div_componentxUDxcentral_parallel_output_13, 
      input_times_b0_div_componentxUDxcentral_parallel_output_14, 
      input_times_b0_div_componentxUDxcentral_parallel_output_15, 
      input_times_b0_div_componentxUDxcentral_parallel_output_16, 
      input_times_b0_div_componentxUDxcentral_parallel_output_17, 
      input_times_b0_div_componentxUDxshifted_substraction_result_0, 
      input_times_b0_mul_componentxUMxFA_127826296_127826240xn3, 
      input_times_b0_mul_componentxUMxFA_127826296_127826240xn2, 
      input_times_b0_mul_componentxUMxAdder_finalxn629, 
      input_times_b0_mul_componentxUMxAdder_finalxn628, 
      input_times_b0_mul_componentxUMxAdder_finalxn607, 
      input_times_b0_mul_componentxUMxAdder_finalxn606, 
      input_times_b0_mul_componentxUMxAdder_finalxn585, 
      input_times_b0_mul_componentxUMxAdder_finalxn584, 
      input_times_b0_mul_componentxUMxAdder_finalxn563, 
      input_times_b0_mul_componentxUMxAdder_finalxn562, 
      input_times_b0_mul_componentxUMxAdder_finalxn541, 
      input_times_b0_mul_componentxUMxAdder_finalxn540, 
      input_times_b0_mul_componentxUMxAdder_finalxn519, 
      input_times_b0_mul_componentxUMxAdder_finalxn518, 
      input_times_b0_mul_componentxUMxAdder_finalxn497, 
      input_times_b0_mul_componentxUMxAdder_finalxn496, 
      input_times_b0_mul_componentxUMxAdder_finalxn475, 
      input_times_b0_mul_componentxUMxAdder_finalxn474, 
      input_times_b0_mul_componentxUMxAdder_finalxn47, 
      input_times_b0_mul_componentxUMxAdder_finalxn25, 
      input_times_b0_mul_componentxUMxAdder_finalxn24, 
      input_times_b0_mul_componentxUMxAdder_finalxn3, 
      input_times_b0_mul_componentxUMxAdder_finalxn2, 
      input_times_b0_div_componentxUDxinput_containerxn40, 
      input_times_b0_div_componentxUDxinput_containerxn38, 
      input_times_b0_div_componentxUDxinput_containerxn37, 
      input_times_b0_div_componentxUDxinput_containerxn36, 
      input_times_b0_div_componentxUDxinput_containerxn35, 
      input_times_b0_div_componentxUDxinput_containerxn34, 
      input_times_b0_div_componentxUDxinput_containerxn33, 
      input_times_b0_div_componentxUDxinput_containerxn32, 
      input_times_b0_div_componentxUDxinput_containerxn31, 
      input_times_b0_div_componentxUDxinput_containerxn30, 
      input_times_b0_div_componentxUDxinput_containerxn29, 
      input_times_b0_div_componentxUDxinput_containerxn28, 
      input_times_b0_div_componentxUDxinput_containerxn27, 
      input_times_b0_div_componentxUDxinput_containerxn26, 
      input_times_b0_div_componentxUDxinput_containerxn25, 
      input_times_b0_div_componentxUDxinput_containerxn24, 
      input_times_b0_div_componentxUDxinput_containerxn23, 
      input_times_b0_div_componentxUDxinput_containerxn22, 
      input_times_b0_div_componentxUDxinput_containerxn21, 
      input_times_b0_div_componentxUDxinput_containerxn20, 
      input_times_b0_div_componentxUDxinput_containerxn19, 
      input_times_b0_div_componentxUDxinput_containerxn18, 
      input_times_b0_div_componentxUDxinput_containerxn17, 
      input_times_b0_div_componentxUDxinput_containerxn16, 
      input_times_b0_div_componentxUDxinput_containerxn15, 
      input_times_b0_div_componentxUDxinput_containerxn14, 
      input_times_b0_div_componentxUDxinput_containerxn13, 
      input_times_b0_div_componentxUDxinput_containerxn12, 
      input_times_b0_div_componentxUDxinput_containerxn11, 
      input_times_b0_div_componentxUDxinput_containerxn10, 
      input_times_b0_div_componentxUDxinput_containerxn9, 
      input_times_b0_div_componentxUDxinput_containerxn8, 
      input_times_b0_div_componentxUDxinput_containerxn7, 
      input_times_b0_div_componentxUDxinput_containerxn6, 
      input_times_b0_div_componentxUDxinput_containerxn5, 
      input_times_b0_div_componentxUDxinput_containerxn3, 
      input_times_b0_div_componentxUDxinput_containerxn2, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_0, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_1, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_2, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_3, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_4, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_5, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_6, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_7, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_8, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_9, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_10, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_11, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_12, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_13, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_14, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_15, 
      input_times_b0_div_componentxUDxinput_containerxparallel_out_16, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn18, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn16, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn14, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn12, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn9, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn8, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn6, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn4, 
      input_times_b0_div_componentxUDxinverter_for_substractionxn2, 
      input_times_b0_div_componentxUDxactually_substractsxn36, 
      input_times_b0_div_componentxUDxactually_substractsxn35, 
      input_times_b0_div_componentxUDxactually_substractsxn34, 
      input_times_b0_div_componentxUDxactually_substractsxn33, 
      input_times_b0_div_componentxUDxactually_substractsxn32, 
      input_times_b0_div_componentxUDxactually_substractsxn31, 
      input_times_b0_div_componentxUDxactually_substractsxn30, 
      input_times_b0_div_componentxUDxactually_substractsxn29, 
      input_times_b0_div_componentxUDxactually_substractsxn28, 
      input_times_b0_div_componentxUDxactually_substractsxn27, 
      input_times_b0_div_componentxUDxactually_substractsxn26, 
      input_times_b0_div_componentxUDxactually_substractsxn25, 
      input_times_b0_div_componentxUDxactually_substractsxn24, 
      input_times_b0_div_componentxUDxactually_substractsxn23, 
      input_times_b0_div_componentxUDxactually_substractsxn18, 
      input_times_b0_div_componentxUDxactually_substractsxn17, 
      input_times_b0_div_componentxUDxactually_substractsxn16, 
      input_times_b0_div_componentxUDxactually_substractsxn15, 
      input_times_b0_div_componentxUDxactually_substractsxn14, 
      input_times_b0_div_componentxUDxactually_substractsxn13, 
      input_times_b0_div_componentxUDxactually_substractsxn12, 
      input_times_b0_div_componentxUDxactually_substractsxn11, 
      input_times_b0_div_componentxUDxactually_substractsxn10, 
      input_times_b0_div_componentxUDxactually_substractsxn9, 
      input_times_b0_div_componentxUDxactually_substractsxn8, 
      input_times_b0_div_componentxUDxactually_substractsxn7, 
      input_times_b0_div_componentxUDxactually_substractsxn6, 
      input_times_b0_div_componentxUDxactually_substractsxn5, 
      input_times_b0_div_componentxUDxactually_substractsxn4, 
      input_times_b0_div_componentxUDxactually_substractsxn3, 
      input_times_b0_div_componentxUDxactually_substractsxn2, 
      input_times_b0_div_componentxUDxactually_substractsxn1, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_1_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_2_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_3_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_4_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_5_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_6_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_7_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_8_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_9_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_10_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_11_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_12_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_13_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_14_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_15_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_16_port, 
      output_p2_times_a2_mul_componentxunsigned_output_inverted_17_port, 
      output_p2_times_a2_mul_componentxunsigned_output_8, 
      output_p2_times_a2_mul_componentxunsigned_output_9, 
      output_p2_times_a2_mul_componentxunsigned_output_10, 
      output_p2_times_a2_mul_componentxunsigned_output_11, 
      output_p2_times_a2_mul_componentxunsigned_output_12, 
      output_p2_times_a2_mul_componentxunsigned_output_13, 
      output_p2_times_a2_mul_componentxunsigned_output_14, 
      output_p2_times_a2_mul_componentxunsigned_output_15, 
      output_p2_times_a2_mul_componentxunsigned_output_16, 
      output_p2_times_a2_mul_componentxunsigned_output_17, 
      output_p2_times_a2_mul_componentxinput_B_inverted_1_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_2_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_3_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_4_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_5_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_6_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_7_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_8_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_9_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_10_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_11_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_12_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_13_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_14_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_15_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_16_port, 
      output_p2_times_a2_mul_componentxinput_B_inverted_17_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_0_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_1_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_2_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_3_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_4_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_5_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_6_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_7_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_8_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_9_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_10_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_11_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_12_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_13_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_14_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_15_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_16_port, 
      output_p2_times_a2_mul_componentxinput_A_inverted_17_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_1_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_2_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_3_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_4_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_5_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_6_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_7_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_8_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_9_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_10_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_11_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_12_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_13_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_14_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_15_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_16_port, 
      output_p1_times_a1_mul_componentxunsigned_output_inverted_17_port, 
      output_p1_times_a1_mul_componentxunsigned_output_8, 
      output_p1_times_a1_mul_componentxunsigned_output_9, 
      output_p1_times_a1_mul_componentxunsigned_output_10, 
      output_p1_times_a1_mul_componentxunsigned_output_11, 
      output_p1_times_a1_mul_componentxunsigned_output_12, 
      output_p1_times_a1_mul_componentxunsigned_output_13, 
      output_p1_times_a1_mul_componentxunsigned_output_14, 
      output_p1_times_a1_mul_componentxunsigned_output_15, 
      output_p1_times_a1_mul_componentxunsigned_output_16, 
      output_p1_times_a1_mul_componentxunsigned_output_17, 
      output_p1_times_a1_mul_componentxinput_B_inverted_1_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_2_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_3_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_4_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_5_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_6_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_7_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_8_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_9_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_10_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_11_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_12_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_13_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_14_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_15_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_16_port, 
      output_p1_times_a1_mul_componentxinput_B_inverted_17_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_0_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_1_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_2_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_3_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_4_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_5_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_6_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_7_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_8_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_9_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_10_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_11_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_12_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_13_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_14_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_15_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_16_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_17_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_1_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_2_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_3_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_4_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_5_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_6_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_7_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_8_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_9_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_10_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_11_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_12_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_13_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_14_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_15_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_16_port, 
      input_p2_times_b2_mul_componentxunsigned_output_inverted_17_port, 
      input_p2_times_b2_mul_componentxunsigned_output_8, 
      input_p2_times_b2_mul_componentxunsigned_output_9, 
      input_p2_times_b2_mul_componentxunsigned_output_10, 
      input_p2_times_b2_mul_componentxunsigned_output_11, 
      input_p2_times_b2_mul_componentxunsigned_output_12, 
      input_p2_times_b2_mul_componentxunsigned_output_13, 
      input_p2_times_b2_mul_componentxunsigned_output_14, 
      input_p2_times_b2_mul_componentxunsigned_output_15, 
      input_p2_times_b2_mul_componentxunsigned_output_16, 
      input_p2_times_b2_mul_componentxunsigned_output_17, 
      input_p2_times_b2_mul_componentxinput_B_inverted_1_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_2_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_3_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_4_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_5_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_6_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_7_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_8_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_9_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_10_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_11_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_12_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_13_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_14_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_15_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_16_port, 
      input_p2_times_b2_mul_componentxinput_B_inverted_17_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_0_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_1_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_2_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_3_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_4_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_5_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_6_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_7_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_8_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_9_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_10_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_11_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_12_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_13_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_14_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_15_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_16_port, 
      input_p2_times_b2_mul_componentxinput_A_inverted_17_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_1_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_2_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_3_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_4_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_5_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_6_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_7_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_8_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_9_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_10_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_11_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_12_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_13_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_14_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_15_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_16_port, 
      input_p1_times_b1_mul_componentxunsigned_output_inverted_17_port, 
      input_p1_times_b1_mul_componentxunsigned_output_8, 
      input_p1_times_b1_mul_componentxunsigned_output_9, 
      input_p1_times_b1_mul_componentxunsigned_output_10, 
      input_p1_times_b1_mul_componentxunsigned_output_11, 
      input_p1_times_b1_mul_componentxunsigned_output_12, 
      input_p1_times_b1_mul_componentxunsigned_output_13, 
      input_p1_times_b1_mul_componentxunsigned_output_14, 
      input_p1_times_b1_mul_componentxunsigned_output_15, 
      input_p1_times_b1_mul_componentxunsigned_output_16, 
      input_p1_times_b1_mul_componentxunsigned_output_17, 
      input_p1_times_b1_mul_componentxinput_B_inverted_1_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_2_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_3_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_4_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_5_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_6_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_7_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_8_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_9_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_10_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_11_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_12_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_13_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_14_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_15_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_16_port, 
      input_p1_times_b1_mul_componentxinput_B_inverted_17_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_0_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_1_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_2_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_3_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_4_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_5_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_6_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_7_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_8_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_9_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_10_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_11_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_12_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_13_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_14_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_15_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_16_port, 
      input_p1_times_b1_mul_componentxinput_A_inverted_17_port, 
      output_p2_times_a2_div_componentxoutput_sign_gated, 
      output_p2_times_a2_div_componentxoutput_sign_gated_prev, 
      output_p2_times_a2_div_componentxunsigned_B_17, 
      output_p2_times_a2_div_componentxunsigned_A_17, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_0_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_1_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_2_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_3_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_4_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_5_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_6_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_7_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_8_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_9_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_10_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_11_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_12_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_13_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_14_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_15_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_16_port, 
      output_p2_times_a2_div_componentxunsigned_output_inverted_17_port, 
      output_p2_times_a2_div_componentxunsigned_output_1, 
      output_p2_times_a2_div_componentxunsigned_output_2, 
      output_p2_times_a2_div_componentxunsigned_output_3, 
      output_p2_times_a2_div_componentxunsigned_output_4, 
      output_p2_times_a2_div_componentxunsigned_output_5, 
      output_p2_times_a2_div_componentxunsigned_output_6, 
      output_p2_times_a2_div_componentxunsigned_output_7, 
      output_p2_times_a2_div_componentxunsigned_output_8, 
      output_p2_times_a2_div_componentxunsigned_output_9, 
      output_p2_times_a2_div_componentxunsigned_output_10, 
      output_p2_times_a2_div_componentxunsigned_output_11, 
      output_p2_times_a2_div_componentxunsigned_output_12, 
      output_p2_times_a2_div_componentxunsigned_output_13, 
      output_p2_times_a2_div_componentxunsigned_output_14, 
      output_p2_times_a2_div_componentxunsigned_output_15, 
      output_p2_times_a2_div_componentxunsigned_output_16, 
      output_p2_times_a2_div_componentxunsigned_output_17, 
      output_p2_times_a2_div_componentxinput_B_inverted_1_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_2_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_3_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_4_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_5_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_6_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_7_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_8_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_9_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_10_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_11_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_12_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_13_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_14_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_15_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_16_port, 
      output_p2_times_a2_div_componentxinput_B_inverted_17_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_1_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_2_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_3_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_4_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_5_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_6_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_7_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_8_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_9_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_10_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_11_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_12_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_13_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_14_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_15_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_16_port, 
      output_p2_times_a2_div_componentxinput_A_inverted_17_port, 
      output_p1_times_a1_div_componentxoutput_sign_gated, 
      output_p1_times_a1_div_componentxoutput_ready_signal, 
      output_p1_times_a1_div_componentxunsigned_B_17, 
      output_p1_times_a1_div_componentxunsigned_A_17, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_0_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_1_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_2_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_3_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_4_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_5_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_6_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_7_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_8_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_9_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_10_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_11_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_12_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_13_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_14_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_15_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_16_port, 
      output_p1_times_a1_div_componentxunsigned_output_inverted_17_port, 
      output_p1_times_a1_div_componentxunsigned_output_1, 
      output_p1_times_a1_div_componentxunsigned_output_2, 
      output_p1_times_a1_div_componentxunsigned_output_3, 
      output_p1_times_a1_div_componentxunsigned_output_4, 
      output_p1_times_a1_div_componentxunsigned_output_5, 
      output_p1_times_a1_div_componentxunsigned_output_6, 
      output_p1_times_a1_div_componentxunsigned_output_7, 
      output_p1_times_a1_div_componentxunsigned_output_8, 
      output_p1_times_a1_div_componentxunsigned_output_9, 
      output_p1_times_a1_div_componentxunsigned_output_10, 
      output_p1_times_a1_div_componentxunsigned_output_11, 
      output_p1_times_a1_div_componentxunsigned_output_12, 
      output_p1_times_a1_div_componentxunsigned_output_13, 
      output_p1_times_a1_div_componentxunsigned_output_14, 
      output_p1_times_a1_div_componentxunsigned_output_15, 
      output_p1_times_a1_div_componentxunsigned_output_16, 
      output_p1_times_a1_div_componentxunsigned_output_17, 
      output_p1_times_a1_div_componentxinput_B_inverted_1_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_2_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_3_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_4_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_5_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_6_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_7_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_8_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_9_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_10_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_11_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_12_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_13_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_14_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_15_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_16_port, 
      output_p1_times_a1_div_componentxinput_B_inverted_17_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_1_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_2_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_3_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_4_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_5_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_6_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_7_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_8_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_9_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_10_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_11_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_12_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_13_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_14_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_15_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_16_port, 
      output_p1_times_a1_div_componentxinput_A_inverted_17_port, 
      input_p2_times_b2_div_componentxoutput_sign_gated, 
      input_p2_times_b2_div_componentxoutput_sign_gated_prev, 
      input_p2_times_b2_div_componentxoutput_ready_signal, 
      input_p2_times_b2_div_componentxunsigned_B_17, 
      input_p2_times_b2_div_componentxunsigned_A_17, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_0_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_1_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_2_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_3_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_4_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_5_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_6_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_7_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_8_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_9_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_10_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_11_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_12_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_13_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_14_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_15_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_16_port, 
      input_p2_times_b2_div_componentxunsigned_output_inverted_17_port, 
      input_p2_times_b2_div_componentxunsigned_output_1, 
      input_p2_times_b2_div_componentxunsigned_output_2, 
      input_p2_times_b2_div_componentxunsigned_output_3, 
      input_p2_times_b2_div_componentxunsigned_output_4, 
      input_p2_times_b2_div_componentxunsigned_output_5, 
      input_p2_times_b2_div_componentxunsigned_output_6, 
      input_p2_times_b2_div_componentxunsigned_output_7, 
      input_p2_times_b2_div_componentxunsigned_output_8, 
      input_p2_times_b2_div_componentxunsigned_output_9, 
      input_p2_times_b2_div_componentxunsigned_output_10, 
      input_p2_times_b2_div_componentxunsigned_output_11, 
      input_p2_times_b2_div_componentxunsigned_output_12, 
      input_p2_times_b2_div_componentxunsigned_output_13, 
      input_p2_times_b2_div_componentxunsigned_output_14, 
      input_p2_times_b2_div_componentxunsigned_output_15, 
      input_p2_times_b2_div_componentxunsigned_output_16, 
      input_p2_times_b2_div_componentxunsigned_output_17, 
      input_p2_times_b2_div_componentxinput_B_inverted_1_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_2_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_3_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_4_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_5_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_6_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_7_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_8_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_9_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_10_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_11_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_12_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_13_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_14_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_15_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_16_port, 
      input_p2_times_b2_div_componentxinput_B_inverted_17_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_1_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_2_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_3_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_4_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_5_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_6_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_7_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_8_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_9_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_10_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_11_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_12_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_13_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_14_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_15_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_16_port, 
      input_p2_times_b2_div_componentxinput_A_inverted_17_port, 
      input_p1_times_b1_div_componentxoutput_sign_gated, 
      input_p1_times_b1_div_componentxoutput_sign_gated_prev, 
      input_p1_times_b1_div_componentxoutput_ready_signal, 
      input_p1_times_b1_div_componentxunsigned_B_17, 
      input_p1_times_b1_div_componentxunsigned_A_17, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_0_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_1_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_2_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_3_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_4_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_5_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_6_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_7_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_8_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_9_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_10_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_11_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_12_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_13_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_14_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_15_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_16_port, 
      input_p1_times_b1_div_componentxunsigned_output_inverted_17_port, 
      input_p1_times_b1_div_componentxunsigned_output_1, 
      input_p1_times_b1_div_componentxunsigned_output_2, 
      input_p1_times_b1_div_componentxunsigned_output_3, 
      input_p1_times_b1_div_componentxunsigned_output_4, 
      input_p1_times_b1_div_componentxunsigned_output_5, 
      input_p1_times_b1_div_componentxunsigned_output_6, 
      input_p1_times_b1_div_componentxunsigned_output_7, 
      input_p1_times_b1_div_componentxunsigned_output_8, 
      input_p1_times_b1_div_componentxunsigned_output_9, 
      input_p1_times_b1_div_componentxunsigned_output_10, 
      input_p1_times_b1_div_componentxunsigned_output_11, 
      input_p1_times_b1_div_componentxunsigned_output_12, 
      input_p1_times_b1_div_componentxunsigned_output_13, 
      input_p1_times_b1_div_componentxunsigned_output_14, 
      input_p1_times_b1_div_componentxunsigned_output_15, 
      input_p1_times_b1_div_componentxunsigned_output_16, 
      input_p1_times_b1_div_componentxunsigned_output_17, 
      input_p1_times_b1_div_componentxinput_B_inverted_1_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_2_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_3_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_4_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_5_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_6_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_7_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_8_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_9_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_10_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_11_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_12_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_13_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_14_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_15_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_16_port, 
      input_p1_times_b1_div_componentxinput_B_inverted_17_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_1_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_2_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_3_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_4_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_5_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_6_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_7_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_8_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_9_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_10_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_11_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_12_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_13_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_14_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_15_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_16_port, 
      input_p1_times_b1_div_componentxinput_A_inverted_17_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_7_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_8_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_9_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_10_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_11_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_12_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_13_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_14_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_15_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_16_port, 
      output_p2_times_a2_mul_componentxUMxsecond_vector_17_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_0_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_1_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_2_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_3_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_4_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_5_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_6_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_7_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_8_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_9_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_10_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_11_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_12_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_13_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_14_port, 
      output_p2_times_a2_mul_componentxUMxfirst_vector_15_port, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128315744_128315968_128316136, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128315464_128315632_128315800, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128220800_128221024_128221136, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128220688_128220856_128220968, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128126256_128220520_128220744, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128125920_128220352_128220576, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128125584_128220184_128220408, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128125248_128219960_128220240, 
      output_p2_times_a2_mul_componentxUMxcarry_layer5_128219792_128220016, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128219792_128220016, 
      output_p2_times_a2_mul_componentxUMxcarry_layer5_128219624_128219848, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128219624_128219848, 
      output_p2_times_a2_mul_componentxUMxcarry_layer5_128219456_128219680, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128219456_128219680, 
      output_p2_times_a2_mul_componentxUMxcarry_layer5_128219288_128219512, 
      output_p2_times_a2_mul_componentxUMxsum_layer5_128219288_128219512, 
      output_p2_times_a2_mul_componentxUMxcarry_layer5_128219120_128219344, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128238312_128238424_128238592, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128237752_128237976_128238144, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128237920_128238088, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128126760_128237640_128237808, 
      output_p2_times_a2_mul_componentxUMxcarry_layer4_128126816_128126928, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128126816_128126928, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128263168_128126424_128126648, 
      output_p2_times_a2_mul_componentxUMxcarry_layer4_128126480_128126592, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128126480_128126592, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128125752_128125976_128126144, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128125416_128125640_128125808, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128125080_128125304_128125472, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128124744_128124968_128125136, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128124632_128124800_128124912, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128247456_128124464_128124688, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128247120_128124240_128124520, 
      output_p2_times_a2_mul_componentxUMxcarry_layer4_128124072_128124296, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128124072_128124296, 
      output_p2_times_a2_mul_componentxUMxcarry_layer4_128123904_128124128, 
      output_p2_times_a2_mul_componentxUMxsum_layer4_128123904_128124128, 
      output_p2_times_a2_mul_componentxUMxcarry_layer4_128123792_128123960, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128264344_128264512, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128263896_128264064_128264176, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128263336_128263560_128263728, 
      output_p2_times_a2_mul_componentxUMxcarry_layer3_128263672_128263840, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128263672_128263840, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128263224_128263392_128263504, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128262664_128262888_128263056, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128262720_128262832_128263000, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128262216_128262384_128262552, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128249696_128249808_128262328, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128197128_128249304_128249528, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128248800_128249024_128249192, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128248296_128248520_128248688, 
      output_p2_times_a2_mul_componentxUMxcarry_layer3_128248464_128248632, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128248464_128248632, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128247960_128248184_128248352, 
      output_p2_times_a2_mul_componentxUMxcarry_layer3_128248016_128248128, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128248016_128248128, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128222880_128247624_128247848, 
      output_p2_times_a2_mul_componentxUMxcarry_layer3_128247680_128247792, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128247680_128247792, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128246952_128247176_128247344, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128246616_128246840_128247008, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128246504_128246672_128246784, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_127827080_128246280_128246560, 
      output_p2_times_a2_mul_componentxUMxcarry_layer3_128246112_128246336, 
      output_p2_times_a2_mul_componentxUMxsum_layer3_128246112_128246336, 
      output_p2_times_a2_mul_componentxUMxcarry_layer3_128246000_128246168, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128199816_128200040_128199984, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128199368_128199480_128199648, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128198864_128199032_128199200, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128198304_128198528_128198696, 
      output_p2_times_a2_mul_componentxUMxcarry_layer2_128198976_128199144, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128198976_128199144, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128198472_128198640_128198808, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128198080_128198192_128198360, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
      output_p2_times_a2_mul_componentxUMxcarry_layer2_128198024_128197968, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128198024_128197968, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128197520_128197632_128197800, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
      output_p2_times_a2_mul_componentxUMxa15_and_b0, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128224952_128225120_128225232, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128224728_128224896_128225064, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128223888_128224112_128224056, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
      output_p2_times_a2_mul_componentxUMxa12_and_b0, 
      output_p2_times_a2_mul_componentxUMxcarry_layer2_128223384_128223552, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128223384_128223552, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128222936_128223104_128223216, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128222376_128222600_128222768, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128222432_128222544_128222712, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128221872_128222096_128222264, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128221760_128221928_128222040, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127635584_128221368_128221592, 
      output_p2_times_a2_mul_componentxUMxa9_and_b0, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127827584_127827808_128221256, 
      output_p2_times_a2_mul_componentxUMxcarry_layer2_127827752_127827920, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127827752_127827920, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127827248_127827472_127827640, 
      output_p2_times_a2_mul_componentxUMxcarry_layer2_127827304_127827416, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127827304_127827416, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
      output_p2_times_a2_mul_componentxUMxa6_and_b0, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127826576_127826800_127826968, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127826464_127826632_127826744, 
      output_p2_times_a2_mul_componentxUMxsum_layer2_127672448_127826240_127826520, 
      output_p2_times_a2_mul_componentxUMxa3_and_b0, 
      output_p2_times_a2_mul_componentxUMxcarry_layer2_127826128_127826296, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127627616_127629520_127824000, 
      output_p2_times_a2_mul_componentxUMxa17_and_b0, 
      output_p2_times_a2_mul_componentxUMxa16_and_b1, 
      output_p2_times_a2_mul_componentxUMxa15_and_b2, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127715984_127849024_127850928, 
      output_p2_times_a2_mul_componentxUMxa14_and_b3, 
      output_p2_times_a2_mul_componentxUMxa13_and_b4, 
      output_p2_times_a2_mul_componentxUMxa12_and_b5, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127636480_127638384_127714080, 
      output_p2_times_a2_mul_componentxUMxa11_and_b6, 
      output_p2_times_a2_mul_componentxUMxa10_and_b7, 
      output_p2_times_a2_mul_componentxUMxa9_and_b8, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127733040_127722720_127724624, 
      output_p2_times_a2_mul_componentxUMxa8_and_b9, 
      output_p2_times_a2_mul_componentxUMxa7_and_b10, 
      output_p2_times_a2_mul_componentxUMxa6_and_b11, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127674016_127675920_127731136, 
      output_p2_times_a2_mul_componentxUMxa5_and_b12, 
      output_p2_times_a2_mul_componentxUMxa4_and_b13, 
      output_p2_times_a2_mul_componentxUMxa3_and_b14, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127832016_127846272_127848176, 
      output_p2_times_a2_mul_componentxUMxa2_and_b15, 
      output_p2_times_a2_mul_componentxUMxa1_and_b16, 
      output_p2_times_a2_mul_componentxUMxa0_and_b17, 
      output_p2_times_a2_mul_componentxUMxcarry_layer1_127627504_127629408, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127627504_127629408, 
      output_p2_times_a2_mul_componentxUMxa16_and_b0, 
      output_p2_times_a2_mul_componentxUMxa15_and_b1, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127715872_127848912_127850816, 
      output_p2_times_a2_mul_componentxUMxa14_and_b2, 
      output_p2_times_a2_mul_componentxUMxa13_and_b3, 
      output_p2_times_a2_mul_componentxUMxa12_and_b4, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127636368_127638272_127713968, 
      output_p2_times_a2_mul_componentxUMxa11_and_b5, 
      output_p2_times_a2_mul_componentxUMxa10_and_b6, 
      output_p2_times_a2_mul_componentxUMxa9_and_b7, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
      output_p2_times_a2_mul_componentxUMxa8_and_b8, 
      output_p2_times_a2_mul_componentxUMxa7_and_b9, 
      output_p2_times_a2_mul_componentxUMxa6_and_b10, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
      output_p2_times_a2_mul_componentxUMxa5_and_b11, 
      output_p2_times_a2_mul_componentxUMxa4_and_b12, 
      output_p2_times_a2_mul_componentxUMxa3_and_b13, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831904_127846160_127848064, 
      output_p2_times_a2_mul_componentxUMxa2_and_b14, 
      output_p2_times_a2_mul_componentxUMxa1_and_b15, 
      output_p2_times_a2_mul_componentxUMxa0_and_b16, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127715760_127848800_127850704, 
      output_p2_times_a2_mul_componentxUMxa14_and_b1, 
      output_p2_times_a2_mul_componentxUMxa13_and_b2, 
      output_p2_times_a2_mul_componentxUMxa12_and_b3, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127636256_127638160_127713856, 
      output_p2_times_a2_mul_componentxUMxa11_and_b4, 
      output_p2_times_a2_mul_componentxUMxa10_and_b5, 
      output_p2_times_a2_mul_componentxUMxa9_and_b6, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732816_127722496_127724400, 
      output_p2_times_a2_mul_componentxUMxa8_and_b7, 
      output_p2_times_a2_mul_componentxUMxa7_and_b8, 
      output_p2_times_a2_mul_componentxUMxa6_and_b9, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
      output_p2_times_a2_mul_componentxUMxa5_and_b10, 
      output_p2_times_a2_mul_componentxUMxa4_and_b11, 
      output_p2_times_a2_mul_componentxUMxa3_and_b12, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
      output_p2_times_a2_mul_componentxUMxa2_and_b13, 
      output_p2_times_a2_mul_componentxUMxa1_and_b14, 
      output_p2_times_a2_mul_componentxUMxa0_and_b15, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
      output_p2_times_a2_mul_componentxUMxa14_and_b0, 
      output_p2_times_a2_mul_componentxUMxa13_and_b1, 
      output_p2_times_a2_mul_componentxUMxa12_and_b2, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127636144_127638048_127713744, 
      output_p2_times_a2_mul_componentxUMxa11_and_b3, 
      output_p2_times_a2_mul_componentxUMxa10_and_b4, 
      output_p2_times_a2_mul_componentxUMxa9_and_b5, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
      output_p2_times_a2_mul_componentxUMxa8_and_b6, 
      output_p2_times_a2_mul_componentxUMxa7_and_b7, 
      output_p2_times_a2_mul_componentxUMxa6_and_b8, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
      output_p2_times_a2_mul_componentxUMxa5_and_b9, 
      output_p2_times_a2_mul_componentxUMxa4_and_b10, 
      output_p2_times_a2_mul_componentxUMxa3_and_b11, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831680_127845936_127847840, 
      output_p2_times_a2_mul_componentxUMxa2_and_b12, 
      output_p2_times_a2_mul_componentxUMxa1_and_b13, 
      output_p2_times_a2_mul_componentxUMxa0_and_b14, 
      output_p2_times_a2_mul_componentxUMxcarry_layer1_127715536_127848576, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127715536_127848576, 
      output_p2_times_a2_mul_componentxUMxa13_and_b0, 
      output_p2_times_a2_mul_componentxUMxa12_and_b1, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
      output_p2_times_a2_mul_componentxUMxa11_and_b2, 
      output_p2_times_a2_mul_componentxUMxa10_and_b3, 
      output_p2_times_a2_mul_componentxUMxa9_and_b4, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
      output_p2_times_a2_mul_componentxUMxa8_and_b5, 
      output_p2_times_a2_mul_componentxUMxa7_and_b6, 
      output_p2_times_a2_mul_componentxUMxa6_and_b7, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673568_127675472_127730688, 
      output_p2_times_a2_mul_componentxUMxa5_and_b8, 
      output_p2_times_a2_mul_componentxUMxa4_and_b9, 
      output_p2_times_a2_mul_componentxUMxa3_and_b10, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
      output_p2_times_a2_mul_componentxUMxa2_and_b11, 
      output_p2_times_a2_mul_componentxUMxa1_and_b12, 
      output_p2_times_a2_mul_componentxUMxa0_and_b13, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127635920_127637824_127713520, 
      output_p2_times_a2_mul_componentxUMxa11_and_b1, 
      output_p2_times_a2_mul_componentxUMxa10_and_b2, 
      output_p2_times_a2_mul_componentxUMxa9_and_b3, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
      output_p2_times_a2_mul_componentxUMxa8_and_b4, 
      output_p2_times_a2_mul_componentxUMxa7_and_b5, 
      output_p2_times_a2_mul_componentxUMxa6_and_b6, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
      output_p2_times_a2_mul_componentxUMxa5_and_b7, 
      output_p2_times_a2_mul_componentxUMxa4_and_b8, 
      output_p2_times_a2_mul_componentxUMxa3_and_b9, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831456_127845712_127847616, 
      output_p2_times_a2_mul_componentxUMxa2_and_b10, 
      output_p2_times_a2_mul_componentxUMxa1_and_b11, 
      output_p2_times_a2_mul_componentxUMxa0_and_b12, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127635808_127637712_127713408, 
      output_p2_times_a2_mul_componentxUMxa11_and_b0, 
      output_p2_times_a2_mul_componentxUMxa10_and_b1, 
      output_p2_times_a2_mul_componentxUMxa9_and_b2, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732368_127722048_127723952, 
      output_p2_times_a2_mul_componentxUMxa8_and_b3, 
      output_p2_times_a2_mul_componentxUMxa7_and_b4, 
      output_p2_times_a2_mul_componentxUMxa6_and_b5, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673344_127675248_127730464, 
      output_p2_times_a2_mul_componentxUMxa5_and_b6, 
      output_p2_times_a2_mul_componentxUMxa4_and_b7, 
      output_p2_times_a2_mul_componentxUMxa3_and_b8, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
      output_p2_times_a2_mul_componentxUMxa2_and_b9, 
      output_p2_times_a2_mul_componentxUMxa1_and_b10, 
      output_p2_times_a2_mul_componentxUMxa0_and_b11, 
      output_p2_times_a2_mul_componentxUMxcarry_layer1_127635696_127637600, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127635696_127637600, 
      output_p2_times_a2_mul_componentxUMxa10_and_b0, 
      output_p2_times_a2_mul_componentxUMxa9_and_b1, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732256_127721936_127723840, 
      output_p2_times_a2_mul_componentxUMxa8_and_b2, 
      output_p2_times_a2_mul_componentxUMxa7_and_b3, 
      output_p2_times_a2_mul_componentxUMxa6_and_b4, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
      output_p2_times_a2_mul_componentxUMxa5_and_b5, 
      output_p2_times_a2_mul_componentxUMxa4_and_b6, 
      output_p2_times_a2_mul_componentxUMxa3_and_b7, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
      output_p2_times_a2_mul_componentxUMxa2_and_b8, 
      output_p2_times_a2_mul_componentxUMxa1_and_b9, 
      output_p2_times_a2_mul_componentxUMxa0_and_b10, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
      output_p2_times_a2_mul_componentxUMxa8_and_b1, 
      output_p2_times_a2_mul_componentxUMxa7_and_b2, 
      output_p2_times_a2_mul_componentxUMxa6_and_b3, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673120_127675024_127730240, 
      output_p2_times_a2_mul_componentxUMxa5_and_b4, 
      output_p2_times_a2_mul_componentxUMxa4_and_b5, 
      output_p2_times_a2_mul_componentxUMxa3_and_b6, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
      output_p2_times_a2_mul_componentxUMxa2_and_b7, 
      output_p2_times_a2_mul_componentxUMxa1_and_b8, 
      output_p2_times_a2_mul_componentxUMxa0_and_b9, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127732032_127721712_127723616, 
      output_p2_times_a2_mul_componentxUMxa8_and_b0, 
      output_p2_times_a2_mul_componentxUMxa7_and_b1, 
      output_p2_times_a2_mul_componentxUMxa6_and_b2, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
      output_p2_times_a2_mul_componentxUMxa5_and_b3, 
      output_p2_times_a2_mul_componentxUMxa4_and_b4, 
      output_p2_times_a2_mul_componentxUMxa3_and_b5, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
      output_p2_times_a2_mul_componentxUMxa2_and_b6, 
      output_p2_times_a2_mul_componentxUMxa1_and_b7, 
      output_p2_times_a2_mul_componentxUMxa0_and_b8, 
      output_p2_times_a2_mul_componentxUMxcarry_layer1_127731920_127721600, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127731920_127721600, 
      output_p2_times_a2_mul_componentxUMxa7_and_b0, 
      output_p2_times_a2_mul_componentxUMxa6_and_b1, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127672896_127674800_127730016, 
      output_p2_times_a2_mul_componentxUMxa5_and_b2, 
      output_p2_times_a2_mul_componentxUMxa4_and_b3, 
      output_p2_times_a2_mul_componentxUMxa3_and_b4, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127830896_127845152_127847056, 
      output_p2_times_a2_mul_componentxUMxa2_and_b5, 
      output_p2_times_a2_mul_componentxUMxa1_and_b6, 
      output_p2_times_a2_mul_componentxUMxa0_and_b7, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127672784_127674688_127729904, 
      output_p2_times_a2_mul_componentxUMxa5_and_b1, 
      output_p2_times_a2_mul_componentxUMxa4_and_b2, 
      output_p2_times_a2_mul_componentxUMxa3_and_b3, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127830784_127845040_127846944, 
      output_p2_times_a2_mul_componentxUMxa2_and_b4, 
      output_p2_times_a2_mul_componentxUMxa1_and_b5, 
      output_p2_times_a2_mul_componentxUMxa0_and_b6, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
      output_p2_times_a2_mul_componentxUMxa5_and_b0, 
      output_p2_times_a2_mul_componentxUMxa4_and_b1, 
      output_p2_times_a2_mul_componentxUMxa3_and_b2, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127830672_127844928_127846832, 
      output_p2_times_a2_mul_componentxUMxa2_and_b3, 
      output_p2_times_a2_mul_componentxUMxa1_and_b4, 
      output_p2_times_a2_mul_componentxUMxa0_and_b5, 
      output_p2_times_a2_mul_componentxUMxcarry_layer1_127672560_127674464, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127672560_127674464, 
      output_p2_times_a2_mul_componentxUMxa4_and_b0, 
      output_p2_times_a2_mul_componentxUMxa3_and_b1, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
      output_p2_times_a2_mul_componentxUMxa2_and_b2, 
      output_p2_times_a2_mul_componentxUMxa1_and_b3, 
      output_p2_times_a2_mul_componentxUMxa0_and_b4, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127830448_127844704_127846608, 
      output_p2_times_a2_mul_componentxUMxa2_and_b1, 
      output_p2_times_a2_mul_componentxUMxa1_and_b2, 
      output_p2_times_a2_mul_componentxUMxa0_and_b3, 
      output_p2_times_a2_mul_componentxUMxsum_layer1_127830336_127844592_127846496, 
      output_p2_times_a2_mul_componentxUMxa2_and_b0, 
      output_p2_times_a2_mul_componentxUMxa1_and_b1, 
      output_p2_times_a2_mul_componentxUMxa0_and_b2, 
      output_p2_times_a2_mul_componentxUMxcarry_layer1_127830168_127844480, 
      output_p2_times_a2_mul_componentxUMxa1_and_b0, 
      output_p2_times_a2_mul_componentxUMxa0_and_b1, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_7_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_8_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_9_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_10_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_11_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_12_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_13_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_14_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_15_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_16_port, 
      output_p1_times_a1_mul_componentxUMxsecond_vector_17_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_0_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_1_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_2_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_3_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_4_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_5_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_6_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_7_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_8_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_9_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_10_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_11_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_12_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_13_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_14_port, 
      output_p1_times_a1_mul_componentxUMxfirst_vector_15_port, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128315744_128315968_128316136, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128315464_128315632_128315800, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128220800_128221024_128221136, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128220688_128220856_128220968, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128126256_128220520_128220744, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128125920_128220352_128220576, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128125584_128220184_128220408, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128125248_128219960_128220240, 
      output_p1_times_a1_mul_componentxUMxcarry_layer5_128219792_128220016, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128219792_128220016, 
      output_p1_times_a1_mul_componentxUMxcarry_layer5_128219624_128219848, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128219624_128219848, 
      output_p1_times_a1_mul_componentxUMxcarry_layer5_128219456_128219680, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128219456_128219680, 
      output_p1_times_a1_mul_componentxUMxcarry_layer5_128219288_128219512, 
      output_p1_times_a1_mul_componentxUMxsum_layer5_128219288_128219512, 
      output_p1_times_a1_mul_componentxUMxcarry_layer5_128219120_128219344, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128238312_128238424_128238592, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128237752_128237976_128238144, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128237920_128238088, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128126760_128237640_128237808, 
      output_p1_times_a1_mul_componentxUMxcarry_layer4_128126816_128126928, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128126816_128126928, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128263168_128126424_128126648, 
      output_p1_times_a1_mul_componentxUMxcarry_layer4_128126480_128126592, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128126480_128126592, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128125752_128125976_128126144, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128125416_128125640_128125808, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128125080_128125304_128125472, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128124744_128124968_128125136, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128124632_128124800_128124912, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128247456_128124464_128124688, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128247120_128124240_128124520, 
      output_p1_times_a1_mul_componentxUMxcarry_layer4_128124072_128124296, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128124072_128124296, 
      output_p1_times_a1_mul_componentxUMxcarry_layer4_128123904_128124128, 
      output_p1_times_a1_mul_componentxUMxsum_layer4_128123904_128124128, 
      output_p1_times_a1_mul_componentxUMxcarry_layer4_128123792_128123960, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128264344_128264512, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128263896_128264064_128264176, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128263336_128263560_128263728, 
      output_p1_times_a1_mul_componentxUMxcarry_layer3_128263672_128263840, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128263672_128263840, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128263224_128263392_128263504, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128262664_128262888_128263056, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128262720_128262832_128263000, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128262216_128262384_128262552, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128249696_128249808_128262328, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128197128_128249304_128249528, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128248800_128249024_128249192, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128248296_128248520_128248688, 
      output_p1_times_a1_mul_componentxUMxcarry_layer3_128248464_128248632, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128248464_128248632, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128247960_128248184_128248352, 
      output_p1_times_a1_mul_componentxUMxcarry_layer3_128248016_128248128, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128248016_128248128, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128222880_128247624_128247848, 
      output_p1_times_a1_mul_componentxUMxcarry_layer3_128247680_128247792, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128247680_128247792, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128246952_128247176_128247344, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128246616_128246840_128247008, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128246504_128246672_128246784, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_127827080_128246280_128246560, 
      output_p1_times_a1_mul_componentxUMxcarry_layer3_128246112_128246336, 
      output_p1_times_a1_mul_componentxUMxsum_layer3_128246112_128246336, 
      output_p1_times_a1_mul_componentxUMxcarry_layer3_128246000_128246168, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128199816_128200040_128199984, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128199368_128199480_128199648, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128198864_128199032_128199200, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128198304_128198528_128198696, 
      output_p1_times_a1_mul_componentxUMxcarry_layer2_128198976_128199144, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128198976_128199144, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128198472_128198640_128198808, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128198080_128198192_128198360, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
      output_p1_times_a1_mul_componentxUMxcarry_layer2_128198024_128197968, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128198024_128197968, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128197520_128197632_128197800, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
      output_p1_times_a1_mul_componentxUMxa15_and_b0, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128224952_128225120_128225232, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128224728_128224896_128225064, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128223888_128224112_128224056, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
      output_p1_times_a1_mul_componentxUMxa12_and_b0, 
      output_p1_times_a1_mul_componentxUMxcarry_layer2_128223384_128223552, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128223384_128223552, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128222936_128223104_128223216, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128222376_128222600_128222768, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128222432_128222544_128222712, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128221872_128222096_128222264, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128221760_128221928_128222040, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127635584_128221368_128221592, 
      output_p1_times_a1_mul_componentxUMxa9_and_b0, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127827584_127827808_128221256, 
      output_p1_times_a1_mul_componentxUMxcarry_layer2_127827752_127827920, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127827752_127827920, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127827248_127827472_127827640, 
      output_p1_times_a1_mul_componentxUMxcarry_layer2_127827304_127827416, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127827304_127827416, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
      output_p1_times_a1_mul_componentxUMxa6_and_b0, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127826576_127826800_127826968, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127826464_127826632_127826744, 
      output_p1_times_a1_mul_componentxUMxsum_layer2_127672448_127826240_127826520, 
      output_p1_times_a1_mul_componentxUMxa3_and_b0, 
      output_p1_times_a1_mul_componentxUMxcarry_layer2_127826128_127826296, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127627616_127629520_127824000, 
      output_p1_times_a1_mul_componentxUMxa17_and_b0, 
      output_p1_times_a1_mul_componentxUMxa16_and_b1, 
      output_p1_times_a1_mul_componentxUMxa15_and_b2, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127715984_127849024_127850928, 
      output_p1_times_a1_mul_componentxUMxa14_and_b3, 
      output_p1_times_a1_mul_componentxUMxa13_and_b4, 
      output_p1_times_a1_mul_componentxUMxa12_and_b5, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127636480_127638384_127714080, 
      output_p1_times_a1_mul_componentxUMxa11_and_b6, 
      output_p1_times_a1_mul_componentxUMxa10_and_b7, 
      output_p1_times_a1_mul_componentxUMxa9_and_b8, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127733040_127722720_127724624, 
      output_p1_times_a1_mul_componentxUMxa8_and_b9, 
      output_p1_times_a1_mul_componentxUMxa7_and_b10, 
      output_p1_times_a1_mul_componentxUMxa6_and_b11, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127674016_127675920_127731136, 
      output_p1_times_a1_mul_componentxUMxa5_and_b12, 
      output_p1_times_a1_mul_componentxUMxa4_and_b13, 
      output_p1_times_a1_mul_componentxUMxa3_and_b14, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127832016_127846272_127848176, 
      output_p1_times_a1_mul_componentxUMxa2_and_b15, 
      output_p1_times_a1_mul_componentxUMxa1_and_b16, 
      output_p1_times_a1_mul_componentxUMxa0_and_b17, 
      output_p1_times_a1_mul_componentxUMxcarry_layer1_127627504_127629408, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127627504_127629408, 
      output_p1_times_a1_mul_componentxUMxa16_and_b0, 
      output_p1_times_a1_mul_componentxUMxa15_and_b1, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127715872_127848912_127850816, 
      output_p1_times_a1_mul_componentxUMxa14_and_b2, 
      output_p1_times_a1_mul_componentxUMxa13_and_b3, 
      output_p1_times_a1_mul_componentxUMxa12_and_b4, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127636368_127638272_127713968, 
      output_p1_times_a1_mul_componentxUMxa11_and_b5, 
      output_p1_times_a1_mul_componentxUMxa10_and_b6, 
      output_p1_times_a1_mul_componentxUMxa9_and_b7, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
      output_p1_times_a1_mul_componentxUMxa8_and_b8, 
      output_p1_times_a1_mul_componentxUMxa7_and_b9, 
      output_p1_times_a1_mul_componentxUMxa6_and_b10, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
      output_p1_times_a1_mul_componentxUMxa5_and_b11, 
      output_p1_times_a1_mul_componentxUMxa4_and_b12, 
      output_p1_times_a1_mul_componentxUMxa3_and_b13, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831904_127846160_127848064, 
      output_p1_times_a1_mul_componentxUMxa2_and_b14, 
      output_p1_times_a1_mul_componentxUMxa1_and_b15, 
      output_p1_times_a1_mul_componentxUMxa0_and_b16, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127715760_127848800_127850704, 
      output_p1_times_a1_mul_componentxUMxa14_and_b1, 
      output_p1_times_a1_mul_componentxUMxa13_and_b2, 
      output_p1_times_a1_mul_componentxUMxa12_and_b3, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127636256_127638160_127713856, 
      output_p1_times_a1_mul_componentxUMxa11_and_b4, 
      output_p1_times_a1_mul_componentxUMxa10_and_b5, 
      output_p1_times_a1_mul_componentxUMxa9_and_b6, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732816_127722496_127724400, 
      output_p1_times_a1_mul_componentxUMxa8_and_b7, 
      output_p1_times_a1_mul_componentxUMxa7_and_b8, 
      output_p1_times_a1_mul_componentxUMxa6_and_b9, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
      output_p1_times_a1_mul_componentxUMxa5_and_b10, 
      output_p1_times_a1_mul_componentxUMxa4_and_b11, 
      output_p1_times_a1_mul_componentxUMxa3_and_b12, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
      output_p1_times_a1_mul_componentxUMxa2_and_b13, 
      output_p1_times_a1_mul_componentxUMxa1_and_b14, 
      output_p1_times_a1_mul_componentxUMxa0_and_b15, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
      output_p1_times_a1_mul_componentxUMxa14_and_b0, 
      output_p1_times_a1_mul_componentxUMxa13_and_b1, 
      output_p1_times_a1_mul_componentxUMxa12_and_b2, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127636144_127638048_127713744, 
      output_p1_times_a1_mul_componentxUMxa11_and_b3, 
      output_p1_times_a1_mul_componentxUMxa10_and_b4, 
      output_p1_times_a1_mul_componentxUMxa9_and_b5, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
      output_p1_times_a1_mul_componentxUMxa8_and_b6, 
      output_p1_times_a1_mul_componentxUMxa7_and_b7, 
      output_p1_times_a1_mul_componentxUMxa6_and_b8, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
      output_p1_times_a1_mul_componentxUMxa5_and_b9, 
      output_p1_times_a1_mul_componentxUMxa4_and_b10, 
      output_p1_times_a1_mul_componentxUMxa3_and_b11, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831680_127845936_127847840, 
      output_p1_times_a1_mul_componentxUMxa2_and_b12, 
      output_p1_times_a1_mul_componentxUMxa1_and_b13, 
      output_p1_times_a1_mul_componentxUMxa0_and_b14, 
      output_p1_times_a1_mul_componentxUMxcarry_layer1_127715536_127848576, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127715536_127848576, 
      output_p1_times_a1_mul_componentxUMxa13_and_b0, 
      output_p1_times_a1_mul_componentxUMxa12_and_b1, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
      output_p1_times_a1_mul_componentxUMxa11_and_b2, 
      output_p1_times_a1_mul_componentxUMxa10_and_b3, 
      output_p1_times_a1_mul_componentxUMxa9_and_b4, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
      output_p1_times_a1_mul_componentxUMxa8_and_b5, 
      output_p1_times_a1_mul_componentxUMxa7_and_b6, 
      output_p1_times_a1_mul_componentxUMxa6_and_b7, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673568_127675472_127730688, 
      output_p1_times_a1_mul_componentxUMxa5_and_b8, 
      output_p1_times_a1_mul_componentxUMxa4_and_b9, 
      output_p1_times_a1_mul_componentxUMxa3_and_b10, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
      output_p1_times_a1_mul_componentxUMxa2_and_b11, 
      output_p1_times_a1_mul_componentxUMxa1_and_b12, 
      output_p1_times_a1_mul_componentxUMxa0_and_b13, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127635920_127637824_127713520, 
      output_p1_times_a1_mul_componentxUMxa11_and_b1, 
      output_p1_times_a1_mul_componentxUMxa10_and_b2, 
      output_p1_times_a1_mul_componentxUMxa9_and_b3, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
      output_p1_times_a1_mul_componentxUMxa8_and_b4, 
      output_p1_times_a1_mul_componentxUMxa7_and_b5, 
      output_p1_times_a1_mul_componentxUMxa6_and_b6, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
      output_p1_times_a1_mul_componentxUMxa5_and_b7, 
      output_p1_times_a1_mul_componentxUMxa4_and_b8, 
      output_p1_times_a1_mul_componentxUMxa3_and_b9, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831456_127845712_127847616, 
      output_p1_times_a1_mul_componentxUMxa2_and_b10, 
      output_p1_times_a1_mul_componentxUMxa1_and_b11, 
      output_p1_times_a1_mul_componentxUMxa0_and_b12, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127635808_127637712_127713408, 
      output_p1_times_a1_mul_componentxUMxa11_and_b0, 
      output_p1_times_a1_mul_componentxUMxa10_and_b1, 
      output_p1_times_a1_mul_componentxUMxa9_and_b2, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732368_127722048_127723952, 
      output_p1_times_a1_mul_componentxUMxa8_and_b3, 
      output_p1_times_a1_mul_componentxUMxa7_and_b4, 
      output_p1_times_a1_mul_componentxUMxa6_and_b5, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673344_127675248_127730464, 
      output_p1_times_a1_mul_componentxUMxa5_and_b6, 
      output_p1_times_a1_mul_componentxUMxa4_and_b7, 
      output_p1_times_a1_mul_componentxUMxa3_and_b8, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
      output_p1_times_a1_mul_componentxUMxa2_and_b9, 
      output_p1_times_a1_mul_componentxUMxa1_and_b10, 
      output_p1_times_a1_mul_componentxUMxa0_and_b11, 
      output_p1_times_a1_mul_componentxUMxcarry_layer1_127635696_127637600, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127635696_127637600, 
      output_p1_times_a1_mul_componentxUMxa10_and_b0, 
      output_p1_times_a1_mul_componentxUMxa9_and_b1, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732256_127721936_127723840, 
      output_p1_times_a1_mul_componentxUMxa8_and_b2, 
      output_p1_times_a1_mul_componentxUMxa7_and_b3, 
      output_p1_times_a1_mul_componentxUMxa6_and_b4, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
      output_p1_times_a1_mul_componentxUMxa5_and_b5, 
      output_p1_times_a1_mul_componentxUMxa4_and_b6, 
      output_p1_times_a1_mul_componentxUMxa3_and_b7, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
      output_p1_times_a1_mul_componentxUMxa2_and_b8, 
      output_p1_times_a1_mul_componentxUMxa1_and_b9, 
      output_p1_times_a1_mul_componentxUMxa0_and_b10, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
      output_p1_times_a1_mul_componentxUMxa8_and_b1, 
      output_p1_times_a1_mul_componentxUMxa7_and_b2, 
      output_p1_times_a1_mul_componentxUMxa6_and_b3, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673120_127675024_127730240, 
      output_p1_times_a1_mul_componentxUMxa5_and_b4, 
      output_p1_times_a1_mul_componentxUMxa4_and_b5, 
      output_p1_times_a1_mul_componentxUMxa3_and_b6, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
      output_p1_times_a1_mul_componentxUMxa2_and_b7, 
      output_p1_times_a1_mul_componentxUMxa1_and_b8, 
      output_p1_times_a1_mul_componentxUMxa0_and_b9, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127732032_127721712_127723616, 
      output_p1_times_a1_mul_componentxUMxa8_and_b0, 
      output_p1_times_a1_mul_componentxUMxa7_and_b1, 
      output_p1_times_a1_mul_componentxUMxa6_and_b2, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
      output_p1_times_a1_mul_componentxUMxa5_and_b3, 
      output_p1_times_a1_mul_componentxUMxa4_and_b4, 
      output_p1_times_a1_mul_componentxUMxa3_and_b5, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
      output_p1_times_a1_mul_componentxUMxa2_and_b6, 
      output_p1_times_a1_mul_componentxUMxa1_and_b7, 
      output_p1_times_a1_mul_componentxUMxa0_and_b8, 
      output_p1_times_a1_mul_componentxUMxcarry_layer1_127731920_127721600, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127731920_127721600, 
      output_p1_times_a1_mul_componentxUMxa7_and_b0, 
      output_p1_times_a1_mul_componentxUMxa6_and_b1, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127672896_127674800_127730016, 
      output_p1_times_a1_mul_componentxUMxa5_and_b2, 
      output_p1_times_a1_mul_componentxUMxa4_and_b3, 
      output_p1_times_a1_mul_componentxUMxa3_and_b4, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127830896_127845152_127847056, 
      output_p1_times_a1_mul_componentxUMxa2_and_b5, 
      output_p1_times_a1_mul_componentxUMxa1_and_b6, 
      output_p1_times_a1_mul_componentxUMxa0_and_b7, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127672784_127674688_127729904, 
      output_p1_times_a1_mul_componentxUMxa5_and_b1, 
      output_p1_times_a1_mul_componentxUMxa4_and_b2, 
      output_p1_times_a1_mul_componentxUMxa3_and_b3, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127830784_127845040_127846944, 
      output_p1_times_a1_mul_componentxUMxa2_and_b4, 
      output_p1_times_a1_mul_componentxUMxa1_and_b5, 
      output_p1_times_a1_mul_componentxUMxa0_and_b6, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
      output_p1_times_a1_mul_componentxUMxa5_and_b0, 
      output_p1_times_a1_mul_componentxUMxa4_and_b1, 
      output_p1_times_a1_mul_componentxUMxa3_and_b2, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127830672_127844928_127846832, 
      output_p1_times_a1_mul_componentxUMxa2_and_b3, 
      output_p1_times_a1_mul_componentxUMxa1_and_b4, 
      output_p1_times_a1_mul_componentxUMxa0_and_b5, 
      output_p1_times_a1_mul_componentxUMxcarry_layer1_127672560_127674464, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127672560_127674464, 
      output_p1_times_a1_mul_componentxUMxa4_and_b0, 
      output_p1_times_a1_mul_componentxUMxa3_and_b1, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
      output_p1_times_a1_mul_componentxUMxa2_and_b2, 
      output_p1_times_a1_mul_componentxUMxa1_and_b3, 
      output_p1_times_a1_mul_componentxUMxa0_and_b4, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127830448_127844704_127846608, 
      output_p1_times_a1_mul_componentxUMxa2_and_b1, 
      output_p1_times_a1_mul_componentxUMxa1_and_b2, 
      output_p1_times_a1_mul_componentxUMxa0_and_b3, 
      output_p1_times_a1_mul_componentxUMxsum_layer1_127830336_127844592_127846496, 
      output_p1_times_a1_mul_componentxUMxa2_and_b0, 
      output_p1_times_a1_mul_componentxUMxa1_and_b1, 
      output_p1_times_a1_mul_componentxUMxa0_and_b2, 
      output_p1_times_a1_mul_componentxUMxcarry_layer1_127830168_127844480, 
      output_p1_times_a1_mul_componentxUMxa1_and_b0, 
      output_p1_times_a1_mul_componentxUMxa0_and_b1, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_7_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_8_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_9_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_10_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_11_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_12_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_13_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_14_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_15_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_16_port, 
      input_p2_times_b2_mul_componentxUMxsecond_vector_17_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_0_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_1_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_2_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_3_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_4_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_5_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_6_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_7_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_8_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_9_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_10_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_11_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_12_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_13_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_14_port, 
      input_p2_times_b2_mul_componentxUMxfirst_vector_15_port, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128315744_128315968_128316136, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128315464_128315632_128315800, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128220800_128221024_128221136, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128220688_128220856_128220968, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128126256_128220520_128220744, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128125920_128220352_128220576, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128125584_128220184_128220408, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128125248_128219960_128220240, 
      input_p2_times_b2_mul_componentxUMxcarry_layer5_128219792_128220016, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128219792_128220016, 
      input_p2_times_b2_mul_componentxUMxcarry_layer5_128219624_128219848, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128219624_128219848, 
      input_p2_times_b2_mul_componentxUMxcarry_layer5_128219456_128219680, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128219456_128219680, 
      input_p2_times_b2_mul_componentxUMxcarry_layer5_128219288_128219512, 
      input_p2_times_b2_mul_componentxUMxsum_layer5_128219288_128219512, 
      input_p2_times_b2_mul_componentxUMxcarry_layer5_128219120_128219344, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128238312_128238424_128238592, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128237752_128237976_128238144, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128237920_128238088, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128126760_128237640_128237808, 
      input_p2_times_b2_mul_componentxUMxcarry_layer4_128126816_128126928, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128126816_128126928, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128263168_128126424_128126648, 
      input_p2_times_b2_mul_componentxUMxcarry_layer4_128126480_128126592, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128126480_128126592, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128125752_128125976_128126144, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128125416_128125640_128125808, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128125080_128125304_128125472, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128124744_128124968_128125136, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128124632_128124800_128124912, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128247456_128124464_128124688, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128247120_128124240_128124520, 
      input_p2_times_b2_mul_componentxUMxcarry_layer4_128124072_128124296, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128124072_128124296, 
      input_p2_times_b2_mul_componentxUMxcarry_layer4_128123904_128124128, 
      input_p2_times_b2_mul_componentxUMxsum_layer4_128123904_128124128, 
      input_p2_times_b2_mul_componentxUMxcarry_layer4_128123792_128123960, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128264344_128264512, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128263896_128264064_128264176, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128263336_128263560_128263728, 
      input_p2_times_b2_mul_componentxUMxcarry_layer3_128263672_128263840, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128263672_128263840, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128263224_128263392_128263504, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128262664_128262888_128263056, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128262720_128262832_128263000, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128262216_128262384_128262552, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128249696_128249808_128262328, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128197128_128249304_128249528, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128248800_128249024_128249192, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128248296_128248520_128248688, 
      input_p2_times_b2_mul_componentxUMxcarry_layer3_128248464_128248632, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128248464_128248632, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128247960_128248184_128248352, 
      input_p2_times_b2_mul_componentxUMxcarry_layer3_128248016_128248128, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128248016_128248128, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128222880_128247624_128247848, 
      input_p2_times_b2_mul_componentxUMxcarry_layer3_128247680_128247792, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128247680_128247792, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128246952_128247176_128247344, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128246616_128246840_128247008, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128246504_128246672_128246784, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_127827080_128246280_128246560, 
      input_p2_times_b2_mul_componentxUMxcarry_layer3_128246112_128246336, 
      input_p2_times_b2_mul_componentxUMxsum_layer3_128246112_128246336, 
      input_p2_times_b2_mul_componentxUMxcarry_layer3_128246000_128246168, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128199816_128200040_128199984, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128199368_128199480_128199648, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128198864_128199032_128199200, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128198304_128198528_128198696, 
      input_p2_times_b2_mul_componentxUMxcarry_layer2_128198976_128199144, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128198976_128199144, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128198472_128198640_128198808, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128198080_128198192_128198360, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
      input_p2_times_b2_mul_componentxUMxcarry_layer2_128198024_128197968, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128198024_128197968, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128197520_128197632_128197800, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
      input_p2_times_b2_mul_componentxUMxa15_and_b0, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128224952_128225120_128225232, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128224728_128224896_128225064, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128223888_128224112_128224056, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
      input_p2_times_b2_mul_componentxUMxa12_and_b0, 
      input_p2_times_b2_mul_componentxUMxcarry_layer2_128223384_128223552, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128223384_128223552, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128222936_128223104_128223216, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128222376_128222600_128222768, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128222432_128222544_128222712, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128221872_128222096_128222264, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128221760_128221928_128222040, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127635584_128221368_128221592, 
      input_p2_times_b2_mul_componentxUMxa9_and_b0, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127827584_127827808_128221256, 
      input_p2_times_b2_mul_componentxUMxcarry_layer2_127827752_127827920, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127827752_127827920, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127827248_127827472_127827640, 
      input_p2_times_b2_mul_componentxUMxcarry_layer2_127827304_127827416, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127827304_127827416, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
      input_p2_times_b2_mul_componentxUMxa6_and_b0, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127826576_127826800_127826968, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127826464_127826632_127826744, 
      input_p2_times_b2_mul_componentxUMxsum_layer2_127672448_127826240_127826520, 
      input_p2_times_b2_mul_componentxUMxa3_and_b0, 
      input_p2_times_b2_mul_componentxUMxcarry_layer2_127826128_127826296, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127627616_127629520_127824000, 
      input_p2_times_b2_mul_componentxUMxa17_and_b0, 
      input_p2_times_b2_mul_componentxUMxa16_and_b1, 
      input_p2_times_b2_mul_componentxUMxa15_and_b2, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127715984_127849024_127850928, 
      input_p2_times_b2_mul_componentxUMxa14_and_b3, 
      input_p2_times_b2_mul_componentxUMxa13_and_b4, 
      input_p2_times_b2_mul_componentxUMxa12_and_b5, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127636480_127638384_127714080, 
      input_p2_times_b2_mul_componentxUMxa11_and_b6, 
      input_p2_times_b2_mul_componentxUMxa10_and_b7, 
      input_p2_times_b2_mul_componentxUMxa9_and_b8, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127733040_127722720_127724624, 
      input_p2_times_b2_mul_componentxUMxa8_and_b9, 
      input_p2_times_b2_mul_componentxUMxa7_and_b10, 
      input_p2_times_b2_mul_componentxUMxa6_and_b11, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127674016_127675920_127731136, 
      input_p2_times_b2_mul_componentxUMxa5_and_b12, 
      input_p2_times_b2_mul_componentxUMxa4_and_b13, 
      input_p2_times_b2_mul_componentxUMxa3_and_b14, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127832016_127846272_127848176, 
      input_p2_times_b2_mul_componentxUMxa2_and_b15, 
      input_p2_times_b2_mul_componentxUMxa1_and_b16, 
      input_p2_times_b2_mul_componentxUMxa0_and_b17, 
      input_p2_times_b2_mul_componentxUMxcarry_layer1_127627504_127629408, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127627504_127629408, 
      input_p2_times_b2_mul_componentxUMxa16_and_b0, 
      input_p2_times_b2_mul_componentxUMxa15_and_b1, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127715872_127848912_127850816, 
      input_p2_times_b2_mul_componentxUMxa14_and_b2, 
      input_p2_times_b2_mul_componentxUMxa13_and_b3, 
      input_p2_times_b2_mul_componentxUMxa12_and_b4, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127636368_127638272_127713968, 
      input_p2_times_b2_mul_componentxUMxa11_and_b5, 
      input_p2_times_b2_mul_componentxUMxa10_and_b6, 
      input_p2_times_b2_mul_componentxUMxa9_and_b7, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
      input_p2_times_b2_mul_componentxUMxa8_and_b8, 
      input_p2_times_b2_mul_componentxUMxa7_and_b9, 
      input_p2_times_b2_mul_componentxUMxa6_and_b10, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
      input_p2_times_b2_mul_componentxUMxa5_and_b11, 
      input_p2_times_b2_mul_componentxUMxa4_and_b12, 
      input_p2_times_b2_mul_componentxUMxa3_and_b13, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831904_127846160_127848064, 
      input_p2_times_b2_mul_componentxUMxa2_and_b14, 
      input_p2_times_b2_mul_componentxUMxa1_and_b15, 
      input_p2_times_b2_mul_componentxUMxa0_and_b16, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127715760_127848800_127850704, 
      input_p2_times_b2_mul_componentxUMxa14_and_b1, 
      input_p2_times_b2_mul_componentxUMxa13_and_b2, 
      input_p2_times_b2_mul_componentxUMxa12_and_b3, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127636256_127638160_127713856, 
      input_p2_times_b2_mul_componentxUMxa11_and_b4, 
      input_p2_times_b2_mul_componentxUMxa10_and_b5, 
      input_p2_times_b2_mul_componentxUMxa9_and_b6, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732816_127722496_127724400, 
      input_p2_times_b2_mul_componentxUMxa8_and_b7, 
      input_p2_times_b2_mul_componentxUMxa7_and_b8, 
      input_p2_times_b2_mul_componentxUMxa6_and_b9, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
      input_p2_times_b2_mul_componentxUMxa5_and_b10, 
      input_p2_times_b2_mul_componentxUMxa4_and_b11, 
      input_p2_times_b2_mul_componentxUMxa3_and_b12, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
      input_p2_times_b2_mul_componentxUMxa2_and_b13, 
      input_p2_times_b2_mul_componentxUMxa1_and_b14, 
      input_p2_times_b2_mul_componentxUMxa0_and_b15, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
      input_p2_times_b2_mul_componentxUMxa14_and_b0, 
      input_p2_times_b2_mul_componentxUMxa13_and_b1, 
      input_p2_times_b2_mul_componentxUMxa12_and_b2, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127636144_127638048_127713744, 
      input_p2_times_b2_mul_componentxUMxa11_and_b3, 
      input_p2_times_b2_mul_componentxUMxa10_and_b4, 
      input_p2_times_b2_mul_componentxUMxa9_and_b5, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
      input_p2_times_b2_mul_componentxUMxa8_and_b6, 
      input_p2_times_b2_mul_componentxUMxa7_and_b7, 
      input_p2_times_b2_mul_componentxUMxa6_and_b8, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
      input_p2_times_b2_mul_componentxUMxa5_and_b9, 
      input_p2_times_b2_mul_componentxUMxa4_and_b10, 
      input_p2_times_b2_mul_componentxUMxa3_and_b11, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831680_127845936_127847840, 
      input_p2_times_b2_mul_componentxUMxa2_and_b12, 
      input_p2_times_b2_mul_componentxUMxa1_and_b13, 
      input_p2_times_b2_mul_componentxUMxa0_and_b14, 
      input_p2_times_b2_mul_componentxUMxcarry_layer1_127715536_127848576, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127715536_127848576, 
      input_p2_times_b2_mul_componentxUMxa13_and_b0, 
      input_p2_times_b2_mul_componentxUMxa12_and_b1, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
      input_p2_times_b2_mul_componentxUMxa11_and_b2, 
      input_p2_times_b2_mul_componentxUMxa10_and_b3, 
      input_p2_times_b2_mul_componentxUMxa9_and_b4, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
      input_p2_times_b2_mul_componentxUMxa8_and_b5, 
      input_p2_times_b2_mul_componentxUMxa7_and_b6, 
      input_p2_times_b2_mul_componentxUMxa6_and_b7, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673568_127675472_127730688, 
      input_p2_times_b2_mul_componentxUMxa5_and_b8, 
      input_p2_times_b2_mul_componentxUMxa4_and_b9, 
      input_p2_times_b2_mul_componentxUMxa3_and_b10, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
      input_p2_times_b2_mul_componentxUMxa2_and_b11, 
      input_p2_times_b2_mul_componentxUMxa1_and_b12, 
      input_p2_times_b2_mul_componentxUMxa0_and_b13, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127635920_127637824_127713520, 
      input_p2_times_b2_mul_componentxUMxa11_and_b1, 
      input_p2_times_b2_mul_componentxUMxa10_and_b2, 
      input_p2_times_b2_mul_componentxUMxa9_and_b3, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
      input_p2_times_b2_mul_componentxUMxa8_and_b4, 
      input_p2_times_b2_mul_componentxUMxa7_and_b5, 
      input_p2_times_b2_mul_componentxUMxa6_and_b6, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
      input_p2_times_b2_mul_componentxUMxa5_and_b7, 
      input_p2_times_b2_mul_componentxUMxa4_and_b8, 
      input_p2_times_b2_mul_componentxUMxa3_and_b9, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831456_127845712_127847616, 
      input_p2_times_b2_mul_componentxUMxa2_and_b10, 
      input_p2_times_b2_mul_componentxUMxa1_and_b11, 
      input_p2_times_b2_mul_componentxUMxa0_and_b12, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127635808_127637712_127713408, 
      input_p2_times_b2_mul_componentxUMxa11_and_b0, 
      input_p2_times_b2_mul_componentxUMxa10_and_b1, 
      input_p2_times_b2_mul_componentxUMxa9_and_b2, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732368_127722048_127723952, 
      input_p2_times_b2_mul_componentxUMxa8_and_b3, 
      input_p2_times_b2_mul_componentxUMxa7_and_b4, 
      input_p2_times_b2_mul_componentxUMxa6_and_b5, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673344_127675248_127730464, 
      input_p2_times_b2_mul_componentxUMxa5_and_b6, 
      input_p2_times_b2_mul_componentxUMxa4_and_b7, 
      input_p2_times_b2_mul_componentxUMxa3_and_b8, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
      input_p2_times_b2_mul_componentxUMxa2_and_b9, 
      input_p2_times_b2_mul_componentxUMxa1_and_b10, 
      input_p2_times_b2_mul_componentxUMxa0_and_b11, 
      input_p2_times_b2_mul_componentxUMxcarry_layer1_127635696_127637600, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127635696_127637600, 
      input_p2_times_b2_mul_componentxUMxa10_and_b0, 
      input_p2_times_b2_mul_componentxUMxa9_and_b1, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732256_127721936_127723840, 
      input_p2_times_b2_mul_componentxUMxa8_and_b2, 
      input_p2_times_b2_mul_componentxUMxa7_and_b3, 
      input_p2_times_b2_mul_componentxUMxa6_and_b4, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
      input_p2_times_b2_mul_componentxUMxa5_and_b5, 
      input_p2_times_b2_mul_componentxUMxa4_and_b6, 
      input_p2_times_b2_mul_componentxUMxa3_and_b7, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
      input_p2_times_b2_mul_componentxUMxa2_and_b8, 
      input_p2_times_b2_mul_componentxUMxa1_and_b9, 
      input_p2_times_b2_mul_componentxUMxa0_and_b10, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
      input_p2_times_b2_mul_componentxUMxa8_and_b1, 
      input_p2_times_b2_mul_componentxUMxa7_and_b2, 
      input_p2_times_b2_mul_componentxUMxa6_and_b3, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673120_127675024_127730240, 
      input_p2_times_b2_mul_componentxUMxa5_and_b4, 
      input_p2_times_b2_mul_componentxUMxa4_and_b5, 
      input_p2_times_b2_mul_componentxUMxa3_and_b6, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
      input_p2_times_b2_mul_componentxUMxa2_and_b7, 
      input_p2_times_b2_mul_componentxUMxa1_and_b8, 
      input_p2_times_b2_mul_componentxUMxa0_and_b9, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127732032_127721712_127723616, 
      input_p2_times_b2_mul_componentxUMxa8_and_b0, 
      input_p2_times_b2_mul_componentxUMxa7_and_b1, 
      input_p2_times_b2_mul_componentxUMxa6_and_b2, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
      input_p2_times_b2_mul_componentxUMxa5_and_b3, 
      input_p2_times_b2_mul_componentxUMxa4_and_b4, 
      input_p2_times_b2_mul_componentxUMxa3_and_b5, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
      input_p2_times_b2_mul_componentxUMxa2_and_b6, 
      input_p2_times_b2_mul_componentxUMxa1_and_b7, 
      input_p2_times_b2_mul_componentxUMxa0_and_b8, 
      input_p2_times_b2_mul_componentxUMxcarry_layer1_127731920_127721600, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127731920_127721600, 
      input_p2_times_b2_mul_componentxUMxa7_and_b0, 
      input_p2_times_b2_mul_componentxUMxa6_and_b1, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127672896_127674800_127730016, 
      input_p2_times_b2_mul_componentxUMxa5_and_b2, 
      input_p2_times_b2_mul_componentxUMxa4_and_b3, 
      input_p2_times_b2_mul_componentxUMxa3_and_b4, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127830896_127845152_127847056, 
      input_p2_times_b2_mul_componentxUMxa2_and_b5, 
      input_p2_times_b2_mul_componentxUMxa1_and_b6, 
      input_p2_times_b2_mul_componentxUMxa0_and_b7, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127672784_127674688_127729904, 
      input_p2_times_b2_mul_componentxUMxa5_and_b1, 
      input_p2_times_b2_mul_componentxUMxa4_and_b2, 
      input_p2_times_b2_mul_componentxUMxa3_and_b3, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127830784_127845040_127846944, 
      input_p2_times_b2_mul_componentxUMxa2_and_b4, 
      input_p2_times_b2_mul_componentxUMxa1_and_b5, 
      input_p2_times_b2_mul_componentxUMxa0_and_b6, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
      input_p2_times_b2_mul_componentxUMxa5_and_b0, 
      input_p2_times_b2_mul_componentxUMxa4_and_b1, 
      input_p2_times_b2_mul_componentxUMxa3_and_b2, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127830672_127844928_127846832, 
      input_p2_times_b2_mul_componentxUMxa2_and_b3, 
      input_p2_times_b2_mul_componentxUMxa1_and_b4, 
      input_p2_times_b2_mul_componentxUMxa0_and_b5, 
      input_p2_times_b2_mul_componentxUMxcarry_layer1_127672560_127674464, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127672560_127674464, 
      input_p2_times_b2_mul_componentxUMxa4_and_b0, 
      input_p2_times_b2_mul_componentxUMxa3_and_b1, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
      input_p2_times_b2_mul_componentxUMxa2_and_b2, 
      input_p2_times_b2_mul_componentxUMxa1_and_b3, 
      input_p2_times_b2_mul_componentxUMxa0_and_b4, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127830448_127844704_127846608, 
      input_p2_times_b2_mul_componentxUMxa2_and_b1, 
      input_p2_times_b2_mul_componentxUMxa1_and_b2, 
      input_p2_times_b2_mul_componentxUMxa0_and_b3, 
      input_p2_times_b2_mul_componentxUMxsum_layer1_127830336_127844592_127846496, 
      input_p2_times_b2_mul_componentxUMxa2_and_b0, 
      input_p2_times_b2_mul_componentxUMxa1_and_b1, 
      input_p2_times_b2_mul_componentxUMxa0_and_b2, 
      input_p2_times_b2_mul_componentxUMxcarry_layer1_127830168_127844480, 
      input_p2_times_b2_mul_componentxUMxa1_and_b0, 
      input_p2_times_b2_mul_componentxUMxa0_and_b1, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_7_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_8_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_9_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_10_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_11_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_12_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_13_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_14_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_15_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_16_port, 
      input_p1_times_b1_mul_componentxUMxsecond_vector_17_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_0_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_1_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_2_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_3_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_4_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_5_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_6_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_7_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_8_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_9_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_10_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_11_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_12_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_13_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_14_port, 
      input_p1_times_b1_mul_componentxUMxfirst_vector_15_port, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128315744_128315968_128316136, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128315464_128315632_128315800, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128220800_128221024_128221136, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128220688_128220856_128220968, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128126256_128220520_128220744, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128125920_128220352_128220576, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128125584_128220184_128220408, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128125248_128219960_128220240, 
      input_p1_times_b1_mul_componentxUMxcarry_layer5_128219792_128220016, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128219792_128220016, 
      input_p1_times_b1_mul_componentxUMxcarry_layer5_128219624_128219848, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128219624_128219848, 
      input_p1_times_b1_mul_componentxUMxcarry_layer5_128219456_128219680, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128219456_128219680, 
      input_p1_times_b1_mul_componentxUMxcarry_layer5_128219288_128219512, 
      input_p1_times_b1_mul_componentxUMxsum_layer5_128219288_128219512, 
      input_p1_times_b1_mul_componentxUMxcarry_layer5_128219120_128219344, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128238312_128238424_128238592, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128237752_128237976_128238144, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128237920_128238088, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128126760_128237640_128237808, 
      input_p1_times_b1_mul_componentxUMxcarry_layer4_128126816_128126928, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128126816_128126928, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128263168_128126424_128126648, 
      input_p1_times_b1_mul_componentxUMxcarry_layer4_128126480_128126592, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128126480_128126592, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128125752_128125976_128126144, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128125416_128125640_128125808, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128125080_128125304_128125472, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128124744_128124968_128125136, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128124632_128124800_128124912, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128247456_128124464_128124688, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128247120_128124240_128124520, 
      input_p1_times_b1_mul_componentxUMxcarry_layer4_128124072_128124296, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128124072_128124296, 
      input_p1_times_b1_mul_componentxUMxcarry_layer4_128123904_128124128, 
      input_p1_times_b1_mul_componentxUMxsum_layer4_128123904_128124128, 
      input_p1_times_b1_mul_componentxUMxcarry_layer4_128123792_128123960, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128264344_128264512, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128263896_128264064_128264176, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128263336_128263560_128263728, 
      input_p1_times_b1_mul_componentxUMxcarry_layer3_128263672_128263840, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128263672_128263840, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128263224_128263392_128263504, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128262664_128262888_128263056, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128262720_128262832_128263000, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128262216_128262384_128262552, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128249696_128249808_128262328, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128197128_128249304_128249528, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128248800_128249024_128249192, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128248296_128248520_128248688, 
      input_p1_times_b1_mul_componentxUMxcarry_layer3_128248464_128248632, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128248464_128248632, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128247960_128248184_128248352, 
      input_p1_times_b1_mul_componentxUMxcarry_layer3_128248016_128248128, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128248016_128248128, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128222880_128247624_128247848, 
      input_p1_times_b1_mul_componentxUMxcarry_layer3_128247680_128247792, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128247680_128247792, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128246952_128247176_128247344, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128246616_128246840_128247008, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128246504_128246672_128246784, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_127827080_128246280_128246560, 
      input_p1_times_b1_mul_componentxUMxcarry_layer3_128246112_128246336, 
      input_p1_times_b1_mul_componentxUMxsum_layer3_128246112_128246336, 
      input_p1_times_b1_mul_componentxUMxcarry_layer3_128246000_128246168, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128199816_128200040_128199984, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128199368_128199480_128199648, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128198864_128199032_128199200, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128198304_128198528_128198696, 
      input_p1_times_b1_mul_componentxUMxcarry_layer2_128198976_128199144, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128198976_128199144, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128198472_128198640_128198808, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128198080_128198192_128198360, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
      input_p1_times_b1_mul_componentxUMxcarry_layer2_128198024_128197968, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128198024_128197968, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128197520_128197632_128197800, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
      input_p1_times_b1_mul_componentxUMxa15_and_b0, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128224952_128225120_128225232, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128224728_128224896_128225064, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128223888_128224112_128224056, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
      input_p1_times_b1_mul_componentxUMxa12_and_b0, 
      input_p1_times_b1_mul_componentxUMxcarry_layer2_128223384_128223552, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128223384_128223552, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128222936_128223104_128223216, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128222376_128222600_128222768, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128222432_128222544_128222712, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128221872_128222096_128222264, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128221760_128221928_128222040, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127635584_128221368_128221592, 
      input_p1_times_b1_mul_componentxUMxa9_and_b0, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127827584_127827808_128221256, 
      input_p1_times_b1_mul_componentxUMxcarry_layer2_127827752_127827920, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127827752_127827920, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127827248_127827472_127827640, 
      input_p1_times_b1_mul_componentxUMxcarry_layer2_127827304_127827416, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127827304_127827416, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
      input_p1_times_b1_mul_componentxUMxa6_and_b0, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127826576_127826800_127826968, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127826464_127826632_127826744, 
      input_p1_times_b1_mul_componentxUMxsum_layer2_127672448_127826240_127826520, 
      input_p1_times_b1_mul_componentxUMxa3_and_b0, 
      input_p1_times_b1_mul_componentxUMxcarry_layer2_127826128_127826296, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127627616_127629520_127824000, 
      input_p1_times_b1_mul_componentxUMxa17_and_b0, 
      input_p1_times_b1_mul_componentxUMxa16_and_b1, 
      input_p1_times_b1_mul_componentxUMxa15_and_b2, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127715984_127849024_127850928, 
      input_p1_times_b1_mul_componentxUMxa14_and_b3, 
      input_p1_times_b1_mul_componentxUMxa13_and_b4, 
      input_p1_times_b1_mul_componentxUMxa12_and_b5, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127636480_127638384_127714080, 
      input_p1_times_b1_mul_componentxUMxa11_and_b6, 
      input_p1_times_b1_mul_componentxUMxa10_and_b7, 
      input_p1_times_b1_mul_componentxUMxa9_and_b8, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127733040_127722720_127724624, 
      input_p1_times_b1_mul_componentxUMxa8_and_b9, 
      input_p1_times_b1_mul_componentxUMxa7_and_b10, 
      input_p1_times_b1_mul_componentxUMxa6_and_b11, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127674016_127675920_127731136, 
      input_p1_times_b1_mul_componentxUMxa5_and_b12, 
      input_p1_times_b1_mul_componentxUMxa4_and_b13, 
      input_p1_times_b1_mul_componentxUMxa3_and_b14, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127832016_127846272_127848176, 
      input_p1_times_b1_mul_componentxUMxa2_and_b15, 
      input_p1_times_b1_mul_componentxUMxa1_and_b16, 
      input_p1_times_b1_mul_componentxUMxa0_and_b17, 
      input_p1_times_b1_mul_componentxUMxcarry_layer1_127627504_127629408, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127627504_127629408, 
      input_p1_times_b1_mul_componentxUMxa16_and_b0, 
      input_p1_times_b1_mul_componentxUMxa15_and_b1, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127715872_127848912_127850816, 
      input_p1_times_b1_mul_componentxUMxa14_and_b2, 
      input_p1_times_b1_mul_componentxUMxa13_and_b3, 
      input_p1_times_b1_mul_componentxUMxa12_and_b4, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127636368_127638272_127713968, 
      input_p1_times_b1_mul_componentxUMxa11_and_b5, 
      input_p1_times_b1_mul_componentxUMxa10_and_b6, 
      input_p1_times_b1_mul_componentxUMxa9_and_b7, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
      input_p1_times_b1_mul_componentxUMxa8_and_b8, 
      input_p1_times_b1_mul_componentxUMxa7_and_b9, 
      input_p1_times_b1_mul_componentxUMxa6_and_b10, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
      input_p1_times_b1_mul_componentxUMxa5_and_b11, 
      input_p1_times_b1_mul_componentxUMxa4_and_b12, 
      input_p1_times_b1_mul_componentxUMxa3_and_b13, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831904_127846160_127848064, 
      input_p1_times_b1_mul_componentxUMxa2_and_b14, 
      input_p1_times_b1_mul_componentxUMxa1_and_b15, 
      input_p1_times_b1_mul_componentxUMxa0_and_b16, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127715760_127848800_127850704, 
      input_p1_times_b1_mul_componentxUMxa14_and_b1, 
      input_p1_times_b1_mul_componentxUMxa13_and_b2, 
      input_p1_times_b1_mul_componentxUMxa12_and_b3, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127636256_127638160_127713856, 
      input_p1_times_b1_mul_componentxUMxa11_and_b4, 
      input_p1_times_b1_mul_componentxUMxa10_and_b5, 
      input_p1_times_b1_mul_componentxUMxa9_and_b6, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732816_127722496_127724400, 
      input_p1_times_b1_mul_componentxUMxa8_and_b7, 
      input_p1_times_b1_mul_componentxUMxa7_and_b8, 
      input_p1_times_b1_mul_componentxUMxa6_and_b9, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
      input_p1_times_b1_mul_componentxUMxa5_and_b10, 
      input_p1_times_b1_mul_componentxUMxa4_and_b11, 
      input_p1_times_b1_mul_componentxUMxa3_and_b12, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
      input_p1_times_b1_mul_componentxUMxa2_and_b13, 
      input_p1_times_b1_mul_componentxUMxa1_and_b14, 
      input_p1_times_b1_mul_componentxUMxa0_and_b15, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
      input_p1_times_b1_mul_componentxUMxa14_and_b0, 
      input_p1_times_b1_mul_componentxUMxa13_and_b1, 
      input_p1_times_b1_mul_componentxUMxa12_and_b2, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127636144_127638048_127713744, 
      input_p1_times_b1_mul_componentxUMxa11_and_b3, 
      input_p1_times_b1_mul_componentxUMxa10_and_b4, 
      input_p1_times_b1_mul_componentxUMxa9_and_b5, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
      input_p1_times_b1_mul_componentxUMxa8_and_b6, 
      input_p1_times_b1_mul_componentxUMxa7_and_b7, 
      input_p1_times_b1_mul_componentxUMxa6_and_b8, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
      input_p1_times_b1_mul_componentxUMxa5_and_b9, 
      input_p1_times_b1_mul_componentxUMxa4_and_b10, 
      input_p1_times_b1_mul_componentxUMxa3_and_b11, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831680_127845936_127847840, 
      input_p1_times_b1_mul_componentxUMxa2_and_b12, 
      input_p1_times_b1_mul_componentxUMxa1_and_b13, 
      input_p1_times_b1_mul_componentxUMxa0_and_b14, 
      input_p1_times_b1_mul_componentxUMxcarry_layer1_127715536_127848576, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127715536_127848576, 
      input_p1_times_b1_mul_componentxUMxa13_and_b0, 
      input_p1_times_b1_mul_componentxUMxa12_and_b1, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
      input_p1_times_b1_mul_componentxUMxa11_and_b2, 
      input_p1_times_b1_mul_componentxUMxa10_and_b3, 
      input_p1_times_b1_mul_componentxUMxa9_and_b4, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
      input_p1_times_b1_mul_componentxUMxa8_and_b5, 
      input_p1_times_b1_mul_componentxUMxa7_and_b6, 
      input_p1_times_b1_mul_componentxUMxa6_and_b7, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673568_127675472_127730688, 
      input_p1_times_b1_mul_componentxUMxa5_and_b8, 
      input_p1_times_b1_mul_componentxUMxa4_and_b9, 
      input_p1_times_b1_mul_componentxUMxa3_and_b10, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
      input_p1_times_b1_mul_componentxUMxa2_and_b11, 
      input_p1_times_b1_mul_componentxUMxa1_and_b12, 
      input_p1_times_b1_mul_componentxUMxa0_and_b13, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127635920_127637824_127713520, 
      input_p1_times_b1_mul_componentxUMxa11_and_b1, 
      input_p1_times_b1_mul_componentxUMxa10_and_b2, 
      input_p1_times_b1_mul_componentxUMxa9_and_b3, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
      input_p1_times_b1_mul_componentxUMxa8_and_b4, 
      input_p1_times_b1_mul_componentxUMxa7_and_b5, 
      input_p1_times_b1_mul_componentxUMxa6_and_b6, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
      input_p1_times_b1_mul_componentxUMxa5_and_b7, 
      input_p1_times_b1_mul_componentxUMxa4_and_b8, 
      input_p1_times_b1_mul_componentxUMxa3_and_b9, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831456_127845712_127847616, 
      input_p1_times_b1_mul_componentxUMxa2_and_b10, 
      input_p1_times_b1_mul_componentxUMxa1_and_b11, 
      input_p1_times_b1_mul_componentxUMxa0_and_b12, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127635808_127637712_127713408, 
      input_p1_times_b1_mul_componentxUMxa11_and_b0, 
      input_p1_times_b1_mul_componentxUMxa10_and_b1, 
      input_p1_times_b1_mul_componentxUMxa9_and_b2, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732368_127722048_127723952, 
      input_p1_times_b1_mul_componentxUMxa8_and_b3, 
      input_p1_times_b1_mul_componentxUMxa7_and_b4, 
      input_p1_times_b1_mul_componentxUMxa6_and_b5, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673344_127675248_127730464, 
      input_p1_times_b1_mul_componentxUMxa5_and_b6, 
      input_p1_times_b1_mul_componentxUMxa4_and_b7, 
      input_p1_times_b1_mul_componentxUMxa3_and_b8, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
      input_p1_times_b1_mul_componentxUMxa2_and_b9, 
      input_p1_times_b1_mul_componentxUMxa1_and_b10, 
      input_p1_times_b1_mul_componentxUMxa0_and_b11, 
      input_p1_times_b1_mul_componentxUMxcarry_layer1_127635696_127637600, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127635696_127637600, 
      input_p1_times_b1_mul_componentxUMxa10_and_b0, 
      input_p1_times_b1_mul_componentxUMxa9_and_b1, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732256_127721936_127723840, 
      input_p1_times_b1_mul_componentxUMxa8_and_b2, 
      input_p1_times_b1_mul_componentxUMxa7_and_b3, 
      input_p1_times_b1_mul_componentxUMxa6_and_b4, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
      input_p1_times_b1_mul_componentxUMxa5_and_b5, 
      input_p1_times_b1_mul_componentxUMxa4_and_b6, 
      input_p1_times_b1_mul_componentxUMxa3_and_b7, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
      input_p1_times_b1_mul_componentxUMxa2_and_b8, 
      input_p1_times_b1_mul_componentxUMxa1_and_b9, 
      input_p1_times_b1_mul_componentxUMxa0_and_b10, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
      input_p1_times_b1_mul_componentxUMxa8_and_b1, 
      input_p1_times_b1_mul_componentxUMxa7_and_b2, 
      input_p1_times_b1_mul_componentxUMxa6_and_b3, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673120_127675024_127730240, 
      input_p1_times_b1_mul_componentxUMxa5_and_b4, 
      input_p1_times_b1_mul_componentxUMxa4_and_b5, 
      input_p1_times_b1_mul_componentxUMxa3_and_b6, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
      input_p1_times_b1_mul_componentxUMxa2_and_b7, 
      input_p1_times_b1_mul_componentxUMxa1_and_b8, 
      input_p1_times_b1_mul_componentxUMxa0_and_b9, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127732032_127721712_127723616, 
      input_p1_times_b1_mul_componentxUMxa8_and_b0, 
      input_p1_times_b1_mul_componentxUMxa7_and_b1, 
      input_p1_times_b1_mul_componentxUMxa6_and_b2, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
      input_p1_times_b1_mul_componentxUMxa5_and_b3, 
      input_p1_times_b1_mul_componentxUMxa4_and_b4, 
      input_p1_times_b1_mul_componentxUMxa3_and_b5, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
      input_p1_times_b1_mul_componentxUMxa2_and_b6, 
      input_p1_times_b1_mul_componentxUMxa1_and_b7, 
      input_p1_times_b1_mul_componentxUMxa0_and_b8, 
      input_p1_times_b1_mul_componentxUMxcarry_layer1_127731920_127721600, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127731920_127721600, 
      input_p1_times_b1_mul_componentxUMxa7_and_b0, 
      input_p1_times_b1_mul_componentxUMxa6_and_b1, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127672896_127674800_127730016, 
      input_p1_times_b1_mul_componentxUMxa5_and_b2, 
      input_p1_times_b1_mul_componentxUMxa4_and_b3, 
      input_p1_times_b1_mul_componentxUMxa3_and_b4, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127830896_127845152_127847056, 
      input_p1_times_b1_mul_componentxUMxa2_and_b5, 
      input_p1_times_b1_mul_componentxUMxa1_and_b6, 
      input_p1_times_b1_mul_componentxUMxa0_and_b7, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127672784_127674688_127729904, 
      input_p1_times_b1_mul_componentxUMxa5_and_b1, 
      input_p1_times_b1_mul_componentxUMxa4_and_b2, 
      input_p1_times_b1_mul_componentxUMxa3_and_b3, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127830784_127845040_127846944, 
      input_p1_times_b1_mul_componentxUMxa2_and_b4, 
      input_p1_times_b1_mul_componentxUMxa1_and_b5, 
      input_p1_times_b1_mul_componentxUMxa0_and_b6, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
      input_p1_times_b1_mul_componentxUMxa5_and_b0, 
      input_p1_times_b1_mul_componentxUMxa4_and_b1, 
      input_p1_times_b1_mul_componentxUMxa3_and_b2, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127830672_127844928_127846832, 
      input_p1_times_b1_mul_componentxUMxa2_and_b3, 
      input_p1_times_b1_mul_componentxUMxa1_and_b4, 
      input_p1_times_b1_mul_componentxUMxa0_and_b5, 
      input_p1_times_b1_mul_componentxUMxcarry_layer1_127672560_127674464, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127672560_127674464, 
      input_p1_times_b1_mul_componentxUMxa4_and_b0, 
      input_p1_times_b1_mul_componentxUMxa3_and_b1, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
      input_p1_times_b1_mul_componentxUMxa2_and_b2, 
      input_p1_times_b1_mul_componentxUMxa1_and_b3, 
      input_p1_times_b1_mul_componentxUMxa0_and_b4, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127830448_127844704_127846608, 
      input_p1_times_b1_mul_componentxUMxa2_and_b1, 
      input_p1_times_b1_mul_componentxUMxa1_and_b2, 
      input_p1_times_b1_mul_componentxUMxa0_and_b3, 
      input_p1_times_b1_mul_componentxUMxsum_layer1_127830336_127844592_127846496, 
      input_p1_times_b1_mul_componentxUMxa2_and_b0, 
      input_p1_times_b1_mul_componentxUMxa1_and_b1, 
      input_p1_times_b1_mul_componentxUMxa0_and_b2, 
      input_p1_times_b1_mul_componentxUMxcarry_layer1_127830168_127844480, 
      input_p1_times_b1_mul_componentxUMxa1_and_b0, 
      input_p1_times_b1_mul_componentxUMxa0_and_b1, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_0_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_1_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_2_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_3_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_4_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_5_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_6_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_7_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_8_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_9_port, 
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_10_port,
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_11_port,
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_12_port,
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_13_port,
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_14_port,
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_15_port,
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_16_port,
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_17_port,
      output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_18_port,
      output_p2_times_a2_div_componentxUDxis_less_than, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_0_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_1_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_2_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_3_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_4_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_5_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_6_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_7_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_8_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_9_port, 
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_10_port,
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_11_port,
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_12_port,
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_13_port,
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_14_port,
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_15_port,
      output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_16_port,
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_1_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_2_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_3_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_4_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_5_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_6_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_7_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_8_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_9_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_10_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_11_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_12_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_13_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_14_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_15_port, 
      output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_16_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_0_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_1_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_2_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_3_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_4_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_5_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_6_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_7_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_8_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_9_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_10_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_11_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_12_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_13_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_14_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_15_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_16_port, 
      output_p2_times_a2_div_componentxUDxquotient_not_gated_17_port, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_0, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_1, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_2, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_3, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_4, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_5, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_6, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_7, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_8, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_9, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_10, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_11, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_12, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_13, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_14, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_15, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_16, 
      output_p2_times_a2_div_componentxUDxcentral_parallel_output_17, 
      output_p2_times_a2_div_componentxUDxshifted_substraction_result_0, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_0_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_1_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_2_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_3_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_4_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_5_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_6_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_7_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_8_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_9_port, 
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_10_port,
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_11_port,
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_12_port,
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_13_port,
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_14_port,
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_15_port,
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_16_port,
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_17_port,
      output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_18_port,
      output_p1_times_a1_div_componentxUDxis_less_than, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_0_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_1_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_2_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_3_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_4_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_5_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_6_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_7_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_8_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_9_port, 
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_10_port,
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_11_port,
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_12_port,
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_13_port,
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_14_port,
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_15_port,
      output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_16_port,
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_1_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_2_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_3_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_4_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_5_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_6_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_7_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_8_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_9_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_10_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_11_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_12_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_13_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_14_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_15_port, 
      output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_16_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_0_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_1_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_2_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_3_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_4_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_5_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_6_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_7_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_8_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_9_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_10_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_11_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_12_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_13_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_14_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_15_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_16_port, 
      output_p1_times_a1_div_componentxUDxquotient_not_gated_17_port, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_0, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_1, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_2, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_3, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_4, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_5, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_6, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_7, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_8, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_9, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_10, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_11, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_12, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_13, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_14, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_15, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_16, 
      output_p1_times_a1_div_componentxUDxcentral_parallel_output_17, 
      output_p1_times_a1_div_componentxUDxshifted_substraction_result_0, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_0_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_1_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_2_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_3_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_4_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_5_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_6_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_7_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_8_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_9_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_10_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_11_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_12_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_13_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_14_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_15_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_16_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_17_port, 
      input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_18_port, 
      input_p2_times_b2_div_componentxUDxis_less_than, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_0_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_1_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_2_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_3_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_4_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_5_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_6_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_7_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_8_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_9_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_10_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_11_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_12_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_13_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_14_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_15_port, 
      input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_16_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_1_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_2_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_3_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_4_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_5_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_6_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_7_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_8_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_9_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_10_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_11_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_12_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_13_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_14_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_15_port, 
      input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_16_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_0_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_1_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_2_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_3_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_4_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_5_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_6_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_7_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_8_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_9_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_10_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_11_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_12_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_13_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_14_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_15_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_16_port, 
      input_p2_times_b2_div_componentxUDxquotient_not_gated_17_port, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_0, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_1, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_2, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_3, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_4, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_5, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_6, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_7, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_8, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_9, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_10, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_11, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_12, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_13, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_14, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_15, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_16, 
      input_p2_times_b2_div_componentxUDxcentral_parallel_output_17, 
      input_p2_times_b2_div_componentxUDxshifted_substraction_result_0, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_0_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_1_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_2_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_3_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_4_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_5_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_6_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_7_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_8_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_9_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_10_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_11_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_12_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_13_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_14_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_15_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_16_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_17_port, 
      input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_18_port, 
      input_p1_times_b1_div_componentxUDxis_less_than, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_0_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_1_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_2_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_3_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_4_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_5_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_6_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_7_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_8_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_9_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_10_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_11_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_12_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_13_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_14_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_15_port, 
      input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_16_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_1_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_2_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_3_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_4_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_5_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_6_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_7_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_8_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_9_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_10_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_11_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_12_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_13_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_14_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_15_port, 
      input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_16_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_0_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_1_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_2_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_3_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_4_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_5_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_6_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_7_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_8_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_9_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_10_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_11_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_12_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_13_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_14_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_15_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_16_port, 
      input_p1_times_b1_div_componentxUDxquotient_not_gated_17_port, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_0, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_1, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_2, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_3, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_4, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_5, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_6, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_7, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_8, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_9, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_10, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_11, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_12, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_13, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_14, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_15, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_16, 
      input_p1_times_b1_div_componentxUDxcentral_parallel_output_17, 
      input_p1_times_b1_div_componentxUDxshifted_substraction_result_0, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_0, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_1, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_2, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_3, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_4, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_5, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_6, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_7, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_8, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_9, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_10, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_11, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_12, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_13, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_14, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_15, 
      output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_16, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_0, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_1, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_2, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_3, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_4, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_5, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_6, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_7, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_8, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_9, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_10, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_11, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_12, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_13, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_14, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_15, 
      output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_16, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_0, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_1, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_2, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_3, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_4, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_5, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_6, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_7, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_8, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_9, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_10, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_11, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_12, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_13, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_14, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_15, 
      input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_16, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_0, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_1, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_2, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_3, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_4, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_5, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_6, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_7, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_8, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_9, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_10, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_11, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_12, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_13, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_14, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_15, 
      input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_16, n1, 
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      change_input_port, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, 
      n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
      n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, 
      n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, 
      n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
      n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
      n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, 
      n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, 
      n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
      n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
      n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
      n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, 
      n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, 
      n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, 
      n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, 
      n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, 
      n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, 
      n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, 
      n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, 
      n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, 
      n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, 
      n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
      n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, 
      n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
      n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, 
      n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, 
      n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, 
      n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, 
      n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
      n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, 
      n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, 
      n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
      n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, 
      n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
      n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, 
      n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, 
      n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, 
      n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, 
      n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, 
      n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, 
      n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, 
      n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
      n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, 
      n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
      n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, 
      n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, 
      n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, 
      n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, 
      n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
      n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
      n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, 
      n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
      n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
      n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
      n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, 
      n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
      n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
      n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
      n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, 
      n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, 
      n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
      n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
      n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, 
      n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, 
      n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
      n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, 
      n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, 
      n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, 
      n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, 
      n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, 
      n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, 
      n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, 
      n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, 
      n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, 
      n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, 
      n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, 
      n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, 
      n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
      n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, 
      n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, 
      n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
      n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
      n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, 
      n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, 
      n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, 
      n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
      n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
      n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
      n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, 
      n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
      n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
      n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, 
      n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, 
      n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, 
      n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
      n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, 
      n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, 
      n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, 
      n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, 
      n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, 
      n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
      n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
      n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
      n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
      n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
      n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
      n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
      n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, 
      n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
      n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, 
      n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
      n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
      n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, 
      n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, 
      n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, 
      n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
      n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
      n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, 
      n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, 
      n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
      n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, 
      n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, 
      n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, 
      n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, 
      n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, 
      n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, 
      n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, 
      n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, 
      n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
      n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, 
      n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, 
      n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
      n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, 
      n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, 
      n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, 
      n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, 
      n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, 
      n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, 
      n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
      n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
      n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, 
      n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, 
      n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, 
      n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, 
      n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, 
      n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, 
      n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
      n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, 
      n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
      n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, 
      n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, 
      n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, 
      n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, 
      n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, 
      n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, 
      n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, 
      n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
      n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, 
      n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
      n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, 
      n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, 
      n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, 
      n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, 
      n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, 
      n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, 
      n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, 
      n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, 
      n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, 
      n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, 
      n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, 
      n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, 
      n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, 
      n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, 
      n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, 
      n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, 
      n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, 
      n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, 
      n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, 
      n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, 
      n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
      n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, 
      n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, 
      n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, 
      n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, 
      n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, 
      n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, 
      n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, 
      n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, 
      n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, 
      n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, 
      n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, 
      n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, 
      n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, 
      n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, 
      n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, 
      n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, 
      n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, 
      n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, 
      n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, 
      n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, 
      n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, 
      n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, 
      n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, 
      n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, 
      n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, 
      n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, 
      n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, 
      n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, 
      n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, 
      n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, 
      n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, 
      n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, 
      n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, 
      n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, 
      n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, 
      n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, 
      n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, 
      n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, 
      n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, 
      n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, 
      n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, 
      n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, 
      n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, 
      n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, 
      n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, 
      n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, 
      n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, 
      n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, 
      n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, 
      n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, 
      n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, 
      n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, 
      n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, 
      n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, 
      n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, 
      n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, 
      n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, 
      n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, 
      n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, 
      n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, 
      n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, 
      n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, 
      n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, 
      n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, 
      n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, 
      n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, 
      n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, 
      n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, 
      n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, 
      n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, 
      n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, 
      n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, 
      n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, 
      n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, 
      n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, 
      n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, 
      n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, 
      n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, 
      n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, 
      n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, 
      n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, 
      n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, 
      n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, 
      n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, 
      n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, 
      n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, 
      n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, 
      n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, 
      n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, 
      n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, 
      n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, 
      n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, 
      n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, 
      n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, 
      n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, 
      n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, 
      n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, 
      n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, 
      n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, 
      n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, 
      n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, 
      n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, 
      n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, 
      n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, 
      n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, 
      n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, 
      n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, 
      n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, 
      n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, 
      n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, 
      n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, 
      n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, 
      n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, 
      n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, 
      n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, 
      n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, 
      n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, 
      n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, 
      n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, 
      n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, 
      n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, 
      n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, 
      n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, 
      n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, 
      n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, 
      n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, 
      n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, 
      n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, 
      n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, 
      n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, 
      n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, 
      n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, 
      n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, 
      n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, 
      n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, 
      n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, 
      n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, 
      n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, 
      n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, 
      n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, 
      n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, 
      n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, 
      n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, 
      n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, 
      n4671, n4672 : std_logic;

begin
   output_signal <= ( output_signal_7_port, output_signal_6_port, 
      output_signal_5_port, output_signal_4_port, output_signal_3_port, 
      output_signal_2_port, output_signal_1_port, 
      output_p1_times_a1_mul_componentxinput_A_inverted_0_port );
   change_input <= change_input_port;
   
   final_adderxU53 : XOR2X4 port map( A => results_a1_a2_inv_0_port, B => 
                           results_b0_b1_b2_0_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_0_port);
   final_adderxU9 : XOR2X4 port map( A => n4166, B => n4167, Y => 
                           output_signal_2_port);
   final_adderxU8 : XOR2X4 port map( A => n4164, B => n4165, Y => 
                           output_signal_3_port);
   final_adderxU7 : XOR2X4 port map( A => n4162, B => n4163, Y => 
                           output_signal_4_port);
   final_adderxU6 : XOR2X4 port map( A => n4160, B => n4161, Y => 
                           output_signal_5_port);
   final_adderxU5 : XOR2X4 port map( A => n4158, B => n4159, Y => 
                           output_signal_6_port);
   final_adderxU4 : XOR2X4 port map( A => n4156, B => n4157, Y => 
                           output_signal_7_port);
   clock_chopper_and_divisionxdivision_ring_reg_1 : DFFSX1 port map( D => 
                           clock_chopper_and_divisionxn47, CK => clk, SN => 
                           n283, Q => 
                           clock_chopper_and_divisionxdivision_ring_1_port, QN 
                           => n1261);
   clock_chopper_and_divisionxdivision_ring_reg_0 : DFFSX1 port map( D => 
                           clock_chopper_and_divisionxn49, CK => clk, SN => 
                           n283, Q => 
                           clock_chopper_and_divisionxdivision_ring_0_port, QN 
                           => n1262);
   clock_chopper_and_divisionxdivision_ring_reg_21 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn26, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_21_port);
   clock_chopper_and_divisionxdivision_ring_reg_20 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn27, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_20_port);
   clock_chopper_and_divisionxdivision_ring_reg_19 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn28, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_19_port);
   clock_chopper_and_divisionxdivision_ring_reg_18 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn29, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_18_port);
   clock_chopper_and_divisionxdivision_ring_reg_17 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn30, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_17_port);
   clock_chopper_and_divisionxdivision_ring_reg_16 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn31, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_16_port);
   clock_chopper_and_divisionxdivision_ring_reg_15 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn32, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_15_port);
   clock_chopper_and_divisionxdivision_ring_reg_14 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn33, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_14_port);
   clock_chopper_and_divisionxdivision_ring_reg_13 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn34, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_13_port);
   clock_chopper_and_divisionxdivision_ring_reg_12 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn35, CK => clk, RN => 
                           n305, Q => 
                           clock_chopper_and_divisionxdivision_ring_12_port);
   clock_chopper_and_divisionxdivision_ring_reg_11 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn36, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_11_port);
   clock_chopper_and_divisionxdivision_ring_reg_10 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn37, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_10_port);
   clock_chopper_and_divisionxdivision_ring_reg_9 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn38, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_9_port);
   clock_chopper_and_divisionxdivision_ring_reg_8 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn39, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_8_port);
   clock_chopper_and_divisionxdivision_ring_reg_7 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn40, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_7_port);
   clock_chopper_and_divisionxdivision_ring_reg_6 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn41, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_6_port);
   clock_chopper_and_divisionxdivision_ring_reg_5 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn42, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_5_port);
   clock_chopper_and_divisionxdivision_ring_reg_4 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn43, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_4_port);
   clock_chopper_and_divisionxdivision_ring_reg_3 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn44, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_3_port);
   clock_chopper_and_divisionxdivision_ring_reg_2 : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn45, CK => clk, RN => 
                           n304, Q => 
                           clock_chopper_and_divisionxdivision_ring_2_port);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn23,
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_16);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn24,
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_15);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn25,
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_14);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn26,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_13);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn27,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_12);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn28,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_11);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn29,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_10);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn30,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_9);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn31,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_8);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn32,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_7);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn33,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_6);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn34,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_5);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn35,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_4);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn36,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_3);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn37,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_2);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn38,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_1);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn40,
                           CK => clk, RN => n301, Q => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_0);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => n2218, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_16);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => n2219, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_15);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => n2220, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_14);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => n2221, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_13);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => n2222, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_12);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => n2223, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_11);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => n2224, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_10);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n2225, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_9);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n2226, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_8);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n2227, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_7);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n2228, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_6);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n2229, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_5);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n2230, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_4);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n2231, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_3);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n2232, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_2);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n2233, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_1);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n2234, CK => clk, RN => n286
                           , Q => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_0);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => n2109, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_16);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => n2110, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_15);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => n2111, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_14);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => n2112, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_13);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => n2113, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_12);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => n2114, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_11);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => n2115, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_10);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n2116, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_9);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n2117, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_8);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n2118, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_7);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n2119, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_6);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n2120, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_5);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n2121, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_4);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n2122, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_3);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n2123, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_2);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n2124, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_1);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n2125, CK => clk, RN => n283
                           , Q => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_0);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => n1999, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_16);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => n2000, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_15);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => n2001, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_14);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => n2002, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_13);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => n2003, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_12);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => n2004, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_11);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => n2005, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_10);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n2006, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_9);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n2007, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_8);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n2008, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_7);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n2009, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_6);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n2010, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_5);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n2011, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_4);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n2012, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_3);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n2013, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_2);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n2014, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_1);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n2015, CK => clk, RN => n295
                           , Q => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_0);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => n1890, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_16);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => n1891, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_15);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => n1892, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_14);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => n1893, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_13);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => n1894, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_12);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => n1895, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_11);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => n1896, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_10);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n1897, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_9);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n1898, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_8);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n1899, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_7);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n1900, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_6);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n1901, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_5);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n1902, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_4);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n1903, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_3);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n1904, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_2);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n1905, CK => clk, RN => n292
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_1);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n1906, CK => clk, RN => n292
                           , Q => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_0);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_19 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_18_port, 
                           CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           );
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_19 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_18_port, 
                           CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxoutput_ready_signal)
                           ;
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_19 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_18_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxoutput_ready_signal)
                           ;
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_17 :
                           DFFRHQX1 port map( D => n2289, CK => clk, RN => n289
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_17_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_17 :
                           DFFRHQX1 port map( D => n2180, CK => clk, RN => n286
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_17_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => n2070, CK => clk, RN => n283
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_17_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => n1961, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_17_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => n1851, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_17_port);
   input_times_b0_div_componentxoutput_sign_gated_prev_reg : DFFRHQX1 port map(
                           D => n379, CK => clk, RN => n305, Q => 
                           input_times_b0_div_componentxoutput_sign_gated_prev)
                           ;
   output_p2_times_a2_div_componentxoutput_sign_gated_prev_reg : DFFRHQX1 port 
                           map( D => n377, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxoutput_sign_gated_prev);
   input_p2_times_b2_div_componentxoutput_sign_gated_prev_reg : DFFRHQX1 port 
                           map( D => n375, CK => clk, RN => n313, Q => 
                           input_p2_times_b2_div_componentxoutput_sign_gated_prev);
   input_p1_times_b1_div_componentxoutput_sign_gated_prev_reg : DFFRHQX1 port 
                           map( D => n373, CK => clk, RN => n313, Q => 
                           input_p1_times_b1_div_componentxoutput_sign_gated_prev);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_16 :
                           DFFRHQX1 port map( D => n2290, CK => clk, RN => n289
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_16_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_15 :
                           DFFRHQX1 port map( D => n2291, CK => clk, RN => n289
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_15_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_14 :
                           DFFRHQX1 port map( D => n2292, CK => clk, RN => n289
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_14_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_13 :
                           DFFRHQX1 port map( D => n2293, CK => clk, RN => n289
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_13_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_12 :
                           DFFRHQX1 port map( D => n2294, CK => clk, RN => n289
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_12_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_11 :
                           DFFRHQX1 port map( D => n2295, CK => clk, RN => n289
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_11_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_10 :
                           DFFRHQX1 port map( D => n2296, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_10_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n2297, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_9_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n2298, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_8_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n2299, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_7_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n2300, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_6_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n2301, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_5_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n2302, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_4_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n2303, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_3_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n2304, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_2_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n2305, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_1_port);
   output_p2_times_a2_div_componentxUDxoutput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n2306, CK => clk, RN => n288
                           , Q => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_0_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_16 :
                           DFFRHQX1 port map( D => n2181, CK => clk, RN => n286
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_16_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_15 :
                           DFFRHQX1 port map( D => n2182, CK => clk, RN => n286
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_15_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_14 :
                           DFFRHQX1 port map( D => n2183, CK => clk, RN => n286
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_14_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_13 :
                           DFFRHQX1 port map( D => n2184, CK => clk, RN => n286
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_13_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_12 :
                           DFFRHQX1 port map( D => n2185, CK => clk, RN => n286
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_12_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_11 :
                           DFFRHQX1 port map( D => n2186, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_11_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_10 :
                           DFFRHQX1 port map( D => n2187, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_10_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n2188, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_9_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n2189, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_8_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n2190, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_7_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n2191, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_6_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n2192, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_5_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n2193, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_4_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n2194, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_3_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n2195, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_2_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n2196, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_1_port);
   output_p1_times_a1_div_componentxUDxoutput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n2197, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_0_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => n2071, CK => clk, RN => n283
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_16_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => n2072, CK => clk, RN => n287
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_15_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => n2073, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_14_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => n2074, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_13_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => n2075, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_12_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => n2076, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_11_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => n2077, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_10_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n2078, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_9_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n2079, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_8_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n2080, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_7_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n2081, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_6_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n2082, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_5_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n2083, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_4_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n2084, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_3_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n2085, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_2_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n2086, CK => clk, RN => n298
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_1_port);
   input_p2_times_b2_div_componentxUDxoutput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n2087, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_0_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => n1962, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_16_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => n1963, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_15_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => n1964, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_14_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => n1965, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_13_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => n1966, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_12_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => n1967, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_11_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => n1968, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_10_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n1969, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_9_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n1970, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_8_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n1971, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_7_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n1972, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_6_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n1973, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_5_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n1974, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_4_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n1975, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_3_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n1976, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_2_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n1977, CK => clk, RN => n295
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_1_port);
   input_p1_times_b1_div_componentxUDxoutput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n1978, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_0_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => n1852, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_16_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => n1853, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_15_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => n1854, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_14_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => n1855, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_13_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => n1856, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_12_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => n1857, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_11_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => n1858, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_10_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n1859, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_9_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n1860, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_8_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n1861, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_7_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n1862, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_6_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n1863, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_5_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n1864, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_4_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n1865, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_3_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n1866, CK => clk, RN => n292
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_2_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n1867, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_1_port);
   input_times_b0_div_componentxUDxoutput_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n1868, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxquotient_not_gated_0_port);
   input_times_b0_div_componentxUDxinput_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxinput_containerxn22,
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxshifted_substraction_result_0);
   output_p2_times_a2_div_componentxUDxinput_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => n2217, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxshifted_substraction_result_0);
   output_p1_times_a1_div_componentxUDxinput_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => n2108, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxshifted_substraction_result_0);
   input_p2_times_b2_div_componentxUDxinput_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => n1998, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxshifted_substraction_result_0);
   input_p1_times_b1_div_componentxUDxinput_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => n1889, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxshifted_substraction_result_0);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_17 
                           : DFFRHQX1 port map( D => n2253, CK => clk, RN => 
                           n288, Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_17);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_17 
                           : DFFRHQX1 port map( D => n2144, CK => clk, RN => 
                           n285, Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_17);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_17 :
                           DFFRHQX1 port map( D => n2034, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_17);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_17 :
                           DFFRHQX1 port map( D => n1925, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_17);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_17 : 
                           DFFRHQX1 port map( D => n1815, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_17);
   clock_chopper_and_divisionxclk_out_reg : DFFRHQX1 port map( D => 
                           clock_chopper_and_divisionxn46, CK => clk, RN => 
                           n304, Q => n4673);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_16 
                           : DFFRHQX1 port map( D => n2254, CK => clk, RN => 
                           n288, Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_16);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_16 
                           : DFFRHQX1 port map( D => n2145, CK => clk, RN => 
                           n285, Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_16);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_16 :
                           DFFRHQX1 port map( D => n2035, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_16);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_16 :
                           DFFRHQX1 port map( D => n1926, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_16);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_16 : 
                           DFFRHQX1 port map( D => n1816, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_16);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_14 
                           : DFFRHQX1 port map( D => n2256, CK => clk, RN => 
                           n288, Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_14);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_14 
                           : DFFRHQX1 port map( D => n2147, CK => clk, RN => 
                           n285, Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_14);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_14 :
                           DFFRHQX1 port map( D => n2037, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_14);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_14 :
                           DFFRHQX1 port map( D => n1928, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_14);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_14 : 
                           DFFRHQX1 port map( D => n1818, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_14);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_15 
                           : DFFRHQX1 port map( D => n2255, CK => clk, RN => 
                           n288, Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_15);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_15 
                           : DFFRHQX1 port map( D => n2146, CK => clk, RN => 
                           n285, Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_15);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_15 :
                           DFFRHQX1 port map( D => n2036, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_15);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_15 :
                           DFFRHQX1 port map( D => n1927, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_15);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_15 : 
                           DFFRHQX1 port map( D => n1817, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_15);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_12 
                           : DFFRHQX1 port map( D => n2258, CK => clk, RN => 
                           n288, Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_12);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_10 
                           : DFFRHQX1 port map( D => n2260, CK => clk, RN => 
                           n287, Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_10);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_8 :
                           DFFRHQX1 port map( D => n2262, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_8);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_12 
                           : DFFRHQX1 port map( D => n2149, CK => clk, RN => 
                           n284, Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_12);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_10 
                           : DFFRHQX1 port map( D => n2151, CK => clk, RN => 
                           n284, Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_10);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_8 :
                           DFFRHQX1 port map( D => n2153, CK => clk, RN => n285
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_8);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_12 :
                           DFFRHQX1 port map( D => n2039, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_12);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_10 :
                           DFFRHQX1 port map( D => n2041, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_10);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n2043, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_8);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_12 :
                           DFFRHQX1 port map( D => n1930, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_12);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_10 :
                           DFFRHQX1 port map( D => n1932, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_10);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n1934, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_8);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_12 : 
                           DFFRHQX1 port map( D => n1820, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_12);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_10 : 
                           DFFRHQX1 port map( D => n1822, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_10);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_8 : 
                           DFFRHQX1 port map( D => n1824, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_8);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_13 
                           : DFFRHQX1 port map( D => n2257, CK => clk, RN => 
                           n288, Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_13);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_11 
                           : DFFRHQX1 port map( D => n2259, CK => clk, RN => 
                           n288, Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_11);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_9 :
                           DFFRHQX1 port map( D => n2261, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_9);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_13 
                           : DFFRHQX1 port map( D => n2148, CK => clk, RN => 
                           n285, Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_13);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_11 
                           : DFFRHQX1 port map( D => n2150, CK => clk, RN => 
                           n284, Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_11);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_9 :
                           DFFRHQX1 port map( D => n2152, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_9);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_13 :
                           DFFRHQX1 port map( D => n2038, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_13);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_11 :
                           DFFRHQX1 port map( D => n2040, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_11);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n2042, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_9);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_13 :
                           DFFRHQX1 port map( D => n1929, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_13);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_11 :
                           DFFRHQX1 port map( D => n1931, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_11);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n1933, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_9);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_13 : 
                           DFFRHQX1 port map( D => n1819, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_13);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_11 : 
                           DFFRHQX1 port map( D => n1821, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_11);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_9 : 
                           DFFRHQX1 port map( D => n1823, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_9);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_6 :
                           DFFRHQX1 port map( D => n2264, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_6);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_4 :
                           DFFRHQX1 port map( D => n2266, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_4);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_6 :
                           DFFRHQX1 port map( D => n2155, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_6);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_4 :
                           DFFRHQX1 port map( D => n2157, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_4);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n2045, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_6);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n2047, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_4);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n1936, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_6);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n1938, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_4);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_6 : 
                           DFFRHQX1 port map( D => n1826, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_6);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_4 : 
                           DFFRHQX1 port map( D => n1828, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_4);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_7 :
                           DFFRHQX1 port map( D => n2263, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_7);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_5 :
                           DFFRHQX1 port map( D => n2265, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_5);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_7 :
                           DFFRHQX1 port map( D => n2154, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_7);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_5 :
                           DFFRHQX1 port map( D => n2156, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_5);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n2044, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_7);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n2046, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_5);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n1935, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_7);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n1937, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_5);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_7 : 
                           DFFRHQX1 port map( D => n1825, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_7);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_5 : 
                           DFFRHQX1 port map( D => n1827, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_5);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_2 :
                           DFFRHQX1 port map( D => n2268, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_2);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_2 :
                           DFFRHQX1 port map( D => n2159, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_2);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n2049, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_2);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n1940, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_2);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_2 : 
                           DFFRHQX1 port map( D => n1830, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_2);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_0 :
                           DFFRHQX1 port map( D => n2270, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_0);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_0 :
                           DFFRHQX1 port map( D => n2161, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_0);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n2051, CK => clk, RN => n296
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_0);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n1942, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_0);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_0 : 
                           DFFRHQX1 port map( D => n1832, CK => clk, RN => n298
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_0);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_1 :
                           DFFRHQX1 port map( D => n2269, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_1);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_1 :
                           DFFRHQX1 port map( D => n2160, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_1);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n2050, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_1);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n1941, CK => clk, RN => n293
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_1);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_1 : 
                           DFFRHQX1 port map( D => n1831, CK => clk, RN => n294
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_1);
   output_p2_times_a2_div_componentxUDxcentral_containerxinternal_value_reg_3 :
                           DFFRHQX1 port map( D => n2267, CK => clk, RN => n287
                           , Q => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_3);
   output_p1_times_a1_div_componentxUDxcentral_containerxinternal_value_reg_3 :
                           DFFRHQX1 port map( D => n2158, CK => clk, RN => n284
                           , Q => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_3);
   input_p2_times_b2_div_componentxUDxcentral_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n2048, CK => clk, RN => n297
                           , Q => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_3);
   input_p1_times_b1_div_componentxUDxcentral_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n1939, CK => clk, RN => n294
                           , Q => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_3);
   input_times_b0_div_componentxUDxcentral_containerxinternal_value_reg_3 : 
                           DFFRHQX1 port map( D => n1829, CK => clk, RN => n291
                           , Q => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_3);
   output_prev_2_registerxq_reg_16 : DFFRHQX1 port map( D => n4671, CK => clk, 
                           RN => n300, Q => output_previous_2_16_port);
   input_prev_2_registerxq_reg_16 : DFFRHQX1 port map( D => n4653, CK => clk, 
                           RN => n299, Q => input_previous_2_16_port);
   output_prev_2_registerxq_reg_14 : DFFRHQX1 port map( D => n4669, CK => clk, 
                           RN => n300, Q => output_previous_2_14_port);
   input_prev_2_registerxq_reg_14 : DFFRHQX1 port map( D => n4651, CK => clk, 
                           RN => n299, Q => input_previous_2_14_port);
   output_prev_2_registerxq_reg_15 : DFFRHQX1 port map( D => n4670, CK => clk, 
                           RN => n300, Q => output_previous_2_15_port);
   input_prev_2_registerxq_reg_15 : DFFRHQX1 port map( D => n4652, CK => clk, 
                           RN => n299, Q => input_previous_2_15_port);
   input_prev_0_registerxq_reg_16 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn18, CK => clk, RN => n305, Q 
                           => input_previous_0_16_port);
   input_prev_1_registerxq_reg_16 : DFFRHQX1 port map( D => n4635, CK => clk, 
                           RN => n313, Q => input_previous_1_16_port);
   input_prev_0_registerxq_reg_15 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn17, CK => clk, RN => n305, Q 
                           => input_previous_0_15_port);
   input_prev_1_registerxq_reg_15 : DFFRHQX1 port map( D => n4634, CK => clk, 
                           RN => n313, Q => input_previous_1_15_port);
   output_prev_2_registerxq_reg_12 : DFFRHQX1 port map( D => n4667, CK => clk, 
                           RN => n300, Q => output_previous_2_12_port);
   input_prev_2_registerxq_reg_12 : DFFRHQX1 port map( D => n4649, CK => clk, 
                           RN => n299, Q => input_previous_2_12_port);
   output_prev_2_registerxq_reg_13 : DFFRHQX1 port map( D => n4668, CK => clk, 
                           RN => n300, Q => output_previous_2_13_port);
   input_prev_2_registerxq_reg_13 : DFFRHQX1 port map( D => n4650, CK => clk, 
                           RN => n299, Q => input_previous_2_13_port);
   input_prev_0_registerxq_reg_14 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn16, CK => clk, RN => n305, Q 
                           => input_previous_0_14_port);
   input_prev_1_registerxq_reg_14 : DFFRHQX1 port map( D => n4633, CK => clk, 
                           RN => n314, Q => input_previous_1_14_port);
   input_prev_0_registerxq_reg_13 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn15, CK => clk, RN => n305, Q 
                           => input_previous_0_13_port);
   input_prev_1_registerxq_reg_13 : DFFRHQX1 port map( D => n4632, CK => clk, 
                           RN => n314, Q => input_previous_1_13_port);
   output_prev_2_registerxq_reg_10 : DFFRHQX1 port map( D => n4665, CK => clk, 
                           RN => n300, Q => output_previous_2_10_port);
   input_prev_2_registerxq_reg_10 : DFFRHQX1 port map( D => n4647, CK => clk, 
                           RN => n299, Q => input_previous_2_10_port);
   output_prev_2_registerxq_reg_11 : DFFRHQX1 port map( D => n4666, CK => clk, 
                           RN => n300, Q => output_previous_2_11_port);
   input_prev_2_registerxq_reg_11 : DFFRHQX1 port map( D => n4648, CK => clk, 
                           RN => n299, Q => input_previous_2_11_port);
   input_prev_0_registerxq_reg_9 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn11, CK => clk, RN => n306, Q 
                           => input_previous_0_9_port);
   output_prev_2_registerxq_reg_9 : DFFRHQX1 port map( D => n4664, CK => clk, 
                           RN => n300, Q => output_previous_2_9_port);
   input_prev_2_registerxq_reg_9 : DFFRHQX1 port map( D => n4646, CK => clk, RN
                           => n299, Q => input_previous_2_9_port);
   input_prev_1_registerxq_reg_9 : DFFRHQX1 port map( D => n4628, CK => clk, RN
                           => n314, Q => input_previous_1_9_port);
   input_prev_0_registerxq_reg_10 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn12, CK => clk, RN => n306, Q 
                           => input_previous_0_10_port);
   input_prev_1_registerxq_reg_10 : DFFRHQX1 port map( D => n4629, CK => clk, 
                           RN => n314, Q => input_previous_1_10_port);
   input_prev_0_registerxq_reg_12 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn14, CK => clk, RN => n305, Q 
                           => input_previous_0_12_port);
   input_prev_1_registerxq_reg_12 : DFFRHQX1 port map( D => n4631, CK => clk, 
                           RN => n314, Q => input_previous_1_12_port);
   input_prev_0_registerxq_reg_11 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn13, CK => clk, RN => n306, Q 
                           => input_previous_0_11_port);
   input_prev_1_registerxq_reg_11 : DFFRHQX1 port map( D => n4630, CK => clk, 
                           RN => n314, Q => input_previous_1_11_port);
   input_prev_0_registerxq_reg_17 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn20, CK => clk, RN => n305, Q 
                           => input_previous_0_17_port);
   output_prev_2_registerxq_reg_17 : DFFRHQX1 port map( D => n4672, CK => clk, 
                           RN => n300, Q => output_previous_2_17_port);
   input_prev_2_registerxq_reg_17 : DFFRHQX1 port map( D => n4654, CK => clk, 
                           RN => n299, Q => input_previous_2_17_port);
   input_prev_1_registerxq_reg_17 : DFFRHQX1 port map( D => n4636, CK => clk, 
                           RN => n313, Q => input_previous_1_17_port);
   output_prev_2_registerxq_reg_4 : DFFRHQX1 port map( D => n4659, CK => clk, 
                           RN => n300, Q => output_previous_2_4_port);
   output_prev_2_registerxq_reg_6 : DFFRHQX1 port map( D => n4661, CK => clk, 
                           RN => n300, Q => output_previous_2_6_port);
   input_prev_2_registerxq_reg_4 : DFFRHQX1 port map( D => n4641, CK => clk, RN
                           => n299, Q => input_previous_2_4_port);
   input_prev_2_registerxq_reg_6 : DFFRHQX1 port map( D => n4643, CK => clk, RN
                           => n299, Q => input_previous_2_6_port);
   output_prev_2_registerxq_reg_8 : DFFRHQX1 port map( D => n4663, CK => clk, 
                           RN => n300, Q => output_previous_2_8_port);
   input_prev_2_registerxq_reg_8 : DFFRHQX1 port map( D => n4645, CK => clk, RN
                           => n299, Q => input_previous_2_8_port);
   output_prev_2_registerxq_reg_3 : DFFRHQX1 port map( D => n4658, CK => clk, 
                           RN => n301, Q => output_previous_2_3_port);
   output_prev_2_registerxq_reg_5 : DFFRHQX1 port map( D => n4660, CK => clk, 
                           RN => n300, Q => output_previous_2_5_port);
   input_prev_2_registerxq_reg_3 : DFFRHQX1 port map( D => n4640, CK => clk, RN
                           => n300, Q => input_previous_2_3_port);
   input_prev_2_registerxq_reg_5 : DFFRHQX1 port map( D => n4642, CK => clk, RN
                           => n299, Q => input_previous_2_5_port);
   output_prev_2_registerxq_reg_7 : DFFRHQX1 port map( D => n4662, CK => clk, 
                           RN => n300, Q => output_previous_2_7_port);
   input_prev_2_registerxq_reg_7 : DFFRHQX1 port map( D => n4644, CK => clk, RN
                           => n299, Q => input_previous_2_7_port);
   input_prev_0_registerxq_reg_4 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn6, CK => clk, RN => n306, Q 
                           => input_previous_0_4_port);
   input_prev_0_registerxq_reg_6 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn8, CK => clk, RN => n306, Q 
                           => input_previous_0_6_port);
   input_prev_1_registerxq_reg_4 : DFFRHQX1 port map( D => n4623, CK => clk, RN
                           => n298, Q => input_previous_1_4_port);
   input_prev_1_registerxq_reg_6 : DFFRHQX1 port map( D => n4625, CK => clk, RN
                           => n298, Q => input_previous_1_6_port);
   input_prev_0_registerxq_reg_8 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn10, CK => clk, RN => n306, Q 
                           => input_previous_0_8_port);
   input_prev_1_registerxq_reg_8 : DFFRHQX1 port map( D => n4627, CK => clk, RN
                           => n314, Q => input_previous_1_8_port);
   input_prev_0_registerxq_reg_3 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn5, CK => clk, RN => n306, Q 
                           => input_previous_0_3_port);
   input_prev_0_registerxq_reg_5 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn7, CK => clk, RN => n306, Q 
                           => input_previous_0_5_port);
   input_prev_1_registerxq_reg_3 : DFFRHQX1 port map( D => n4622, CK => clk, RN
                           => n299, Q => input_previous_1_3_port);
   input_prev_1_registerxq_reg_5 : DFFRHQX1 port map( D => n4624, CK => clk, RN
                           => n298, Q => input_previous_1_5_port);
   input_prev_0_registerxq_reg_7 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn9, CK => clk, RN => n306, Q 
                           => input_previous_0_7_port);
   input_prev_1_registerxq_reg_7 : DFFRHQX1 port map( D => n4626, CK => clk, RN
                           => n302, Q => input_previous_1_7_port);
   output_prev_2_registerxq_reg_2 : DFFRHQX1 port map( D => n4657, CK => clk, 
                           RN => n301, Q => output_previous_2_2_port);
   input_prev_2_registerxq_reg_2 : DFFRHQX1 port map( D => n4639, CK => clk, RN
                           => n300, Q => input_previous_2_2_port);
   output_prev_2_registerxq_reg_1 : DFFRHQX1 port map( D => n4656, CK => clk, 
                           RN => n301, Q => output_previous_2_1_port);
   input_prev_2_registerxq_reg_1 : DFFRHQX1 port map( D => n4638, CK => clk, RN
                           => n300, Q => input_previous_2_1_port);
   input_prev_0_registerxq_reg_2 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn4, CK => clk, RN => n306, Q 
                           => input_previous_0_2_port);
   input_prev_1_registerxq_reg_2 : DFFRHQX1 port map( D => n4621, CK => clk, RN
                           => n299, Q => input_previous_1_2_port);
   input_prev_0_registerxq_reg_1 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn3, CK => clk, RN => n306, Q 
                           => input_previous_0_1_port);
   input_prev_1_registerxq_reg_1 : DFFRHQX1 port map( D => n4620, CK => clk, RN
                           => n299, Q => input_previous_1_1_port);
   output_prev_2_registerxq_reg_0 : DFFRHQX1 port map( D => n4655, CK => clk, 
                           RN => n301, Q => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_0_port);
   input_prev_2_registerxq_reg_0 : DFFRHQX1 port map( D => n4637, CK => clk, RN
                           => n300, Q => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_0_port);
   input_prev_0_registerxq_reg_0 : DFFRHQX1 port map( D => 
                           input_prev_0_registerxn2, CK => clk, RN => n283, Q 
                           => 
                           input_times_b0_mul_componentxinput_A_inverted_0_port
                           );
   input_prev_1_registerxq_reg_0 : DFFRHQX1 port map( D => n4619, CK => clk, RN
                           => n299, Q => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_0_port);
   input_times_b0_div_componentxUDxquotient_reg_17 : DFFRHQX1 port map( D => 
                           n1281, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_17);
   output_p2_times_a2_div_componentxUDxquotient_reg_17 : DFFRHQX1 port map( D 
                           => n1400, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_17)
                           ;
   output_p1_times_a1_div_componentxUDxquotient_reg_17 : DFFRHQX1 port map( D 
                           => n1419, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_17)
                           ;
   input_p2_times_b2_div_componentxUDxquotient_reg_17 : DFFRHQX1 port map( D =>
                           n1438, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_17);
   input_p1_times_b1_div_componentxUDxquotient_reg_17 : DFFRHQX1 port map( D =>
                           n1457, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_17);
   output_p2_times_a2_div_componentxUDxquotient_reg_16 : DFFRHQX1 port map( D 
                           => n1399, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_16)
                           ;
   output_p1_times_a1_div_componentxUDxquotient_reg_16 : DFFRHQX1 port map( D 
                           => n1418, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_16)
                           ;
   input_p2_times_b2_div_componentxUDxquotient_reg_16 : DFFRHQX1 port map( D =>
                           n1437, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_16);
   input_times_b0_div_componentxUDxquotient_reg_16 : DFFRHQX1 port map( D => 
                           n1280, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_16);
   input_p1_times_b1_div_componentxUDxquotient_reg_16 : DFFRHQX1 port map( D =>
                           n1456, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_16);
   input_p2_times_b2_div_componentxUDxquotient_reg_12 : DFFRHQX1 port map( D =>
                           n1433, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_12);
   input_times_b0_div_componentxUDxquotient_reg_14 : DFFRHQX1 port map( D => 
                           n1278, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_14);
   output_p2_times_a2_div_componentxUDxquotient_reg_14 : DFFRHQX1 port map( D 
                           => n1397, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_14)
                           ;
   output_p1_times_a1_div_componentxUDxquotient_reg_14 : DFFRHQX1 port map( D 
                           => n1416, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_14)
                           ;
   input_p2_times_b2_div_componentxUDxquotient_reg_14 : DFFRHQX1 port map( D =>
                           n1435, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_14);
   input_p1_times_b1_div_componentxUDxquotient_reg_14 : DFFRHQX1 port map( D =>
                           n1454, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_14);
   input_times_b0_div_componentxUDxquotient_reg_15 : DFFRHQX1 port map( D => 
                           n1279, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_15);
   output_p2_times_a2_div_componentxUDxquotient_reg_15 : DFFRHQX1 port map( D 
                           => n1398, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_15)
                           ;
   output_p1_times_a1_div_componentxUDxquotient_reg_15 : DFFRHQX1 port map( D 
                           => n1417, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_15)
                           ;
   input_p2_times_b2_div_componentxUDxquotient_reg_15 : DFFRHQX1 port map( D =>
                           n1436, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_15);
   input_p1_times_b1_div_componentxUDxquotient_reg_15 : DFFRHQX1 port map( D =>
                           n1455, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_15);
   input_p2_times_b2_div_componentxUDxquotient_reg_11 : DFFRHQX1 port map( D =>
                           n1432, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_11);
   output_p1_times_a1_div_componentxUDxquotient_reg_13 : DFFRHQX1 port map( D 
                           => n1415, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_13)
                           ;
   input_p2_times_b2_div_componentxUDxquotient_reg_13 : DFFRHQX1 port map( D =>
                           n1434, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_13);
   input_times_b0_div_componentxUDxquotient_reg_10 : DFFRHQX1 port map( D => 
                           n1274, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_10);
   output_p2_times_a2_div_componentxUDxquotient_reg_10 : DFFRHQX1 port map( D 
                           => n1393, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_10)
                           ;
   output_p1_times_a1_div_componentxUDxquotient_reg_10 : DFFRHQX1 port map( D 
                           => n1412, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_10)
                           ;
   input_p2_times_b2_div_componentxUDxquotient_reg_10 : DFFRHQX1 port map( D =>
                           n1431, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_10);
   input_p1_times_b1_div_componentxUDxquotient_reg_10 : DFFRHQX1 port map( D =>
                           n1450, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_10);
   input_times_b0_div_componentxUDxquotient_reg_12 : DFFRHQX1 port map( D => 
                           n1276, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_12);
   output_p2_times_a2_div_componentxUDxquotient_reg_12 : DFFRHQX1 port map( D 
                           => n1395, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_12)
                           ;
   output_p1_times_a1_div_componentxUDxquotient_reg_12 : DFFRHQX1 port map( D 
                           => n1414, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_12)
                           ;
   input_p1_times_b1_div_componentxUDxquotient_reg_12 : DFFRHQX1 port map( D =>
                           n1452, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_12);
   input_p2_times_b2_div_componentxUDxquotient_reg_8 : DFFRHQX1 port map( D => 
                           n1428, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_8);
   input_times_b0_div_componentxUDxquotient_reg_11 : DFFRHQX1 port map( D => 
                           n1275, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_11);
   output_p2_times_a2_div_componentxUDxquotient_reg_11 : DFFRHQX1 port map( D 
                           => n1394, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_11)
                           ;
   output_p1_times_a1_div_componentxUDxquotient_reg_11 : DFFRHQX1 port map( D 
                           => n1413, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_11)
                           ;
   input_p1_times_b1_div_componentxUDxquotient_reg_11 : DFFRHQX1 port map( D =>
                           n1451, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_11);
   input_times_b0_div_componentxUDxquotient_reg_9 : DFFRHQX1 port map( D => 
                           n1273, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_9);
   output_p2_times_a2_div_componentxUDxquotient_reg_9 : DFFRHQX1 port map( D =>
                           n1392, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_9);
   output_p1_times_a1_div_componentxUDxquotient_reg_9 : DFFRHQX1 port map( D =>
                           n1411, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_9);
   input_p2_times_b2_div_componentxUDxquotient_reg_9 : DFFRHQX1 port map( D => 
                           n1430, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_9);
   input_times_b0_div_componentxUDxquotient_reg_13 : DFFRHQX1 port map( D => 
                           n1277, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_13);
   output_p2_times_a2_div_componentxUDxquotient_reg_13 : DFFRHQX1 port map( D 
                           => n1396, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_13)
                           ;
   input_p2_times_b2_div_componentxUDxquotient_reg_7 : DFFRHQX1 port map( D => 
                           n1427, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_7);
   input_p1_times_b1_div_componentxUDxquotient_reg_13 : DFFRHQX1 port map( D =>
                           n1453, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_13);
   input_p2_times_b2_div_componentxUDxquotient_reg_2 : DFFRHQX1 port map( D => 
                           n1422, CK => clk, RN => n309, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_2);
   input_times_b0_div_componentxUDxquotient_reg_6 : DFFRHQX1 port map( D => 
                           n1269, CK => clk, RN => n304, Q => 
                           input_times_b0_div_componentxunsigned_output_6);
   output_p2_times_a2_div_componentxUDxquotient_reg_6 : DFFRHQX1 port map( D =>
                           n1388, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_6);
   output_p1_times_a1_div_componentxUDxquotient_reg_6 : DFFRHQX1 port map( D =>
                           n1407, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_6);
   input_p2_times_b2_div_componentxUDxquotient_reg_4 : DFFRHQX1 port map( D => 
                           n1424, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_4);
   input_p2_times_b2_div_componentxUDxquotient_reg_6 : DFFRHQX1 port map( D => 
                           n1426, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_6);
   input_p1_times_b1_div_componentxUDxquotient_reg_6 : DFFRHQX1 port map( D => 
                           n1445, CK => clk, RN => n306, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_6);
   input_times_b0_div_componentxUDxquotient_reg_8 : DFFRHQX1 port map( D => 
                           n1271, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_8);
   output_p2_times_a2_div_componentxUDxquotient_reg_8 : DFFRHQX1 port map( D =>
                           n1390, CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_8);
   output_p1_times_a1_div_componentxUDxquotient_reg_8 : DFFRHQX1 port map( D =>
                           n1409, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_8);
   input_p1_times_b1_div_componentxUDxquotient_reg_8 : DFFRHQX1 port map( D => 
                           n1447, CK => clk, RN => n310, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_8);
   input_times_b0_div_componentxUDxquotient_reg_5 : DFFRHQX1 port map( D => 
                           n1268, CK => clk, RN => n304, Q => 
                           input_times_b0_div_componentxunsigned_output_5);
   output_p2_times_a2_div_componentxUDxquotient_reg_5 : DFFRHQX1 port map( D =>
                           n1387, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_5);
   output_p1_times_a1_div_componentxUDxquotient_reg_5 : DFFRHQX1 port map( D =>
                           n1406, CK => clk, RN => n311, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_5);
   input_p2_times_b2_div_componentxUDxquotient_reg_3 : DFFRHQX1 port map( D => 
                           n1423, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_3);
   input_p2_times_b2_div_componentxUDxquotient_reg_5 : DFFRHQX1 port map( D => 
                           n1425, CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_5);
   input_p1_times_b1_div_componentxUDxquotient_reg_5 : DFFRHQX1 port map( D => 
                           n1444, CK => clk, RN => n306, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_5);
   input_p1_times_b1_div_componentxUDxquotient_reg_9 : DFFRHQX1 port map( D => 
                           n1449, CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_9);
   input_times_b0_div_componentxUDxquotient_reg_7 : DFFRHQX1 port map( D => 
                           n1270, CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxunsigned_output_7);
   output_p2_times_a2_div_componentxUDxquotient_reg_7 : DFFRHQX1 port map( D =>
                           n1389, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_7);
   output_p1_times_a1_div_componentxUDxquotient_reg_7 : DFFRHQX1 port map( D =>
                           n1408, CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_7);
   input_p1_times_b1_div_componentxUDxquotient_reg_7 : DFFRHQX1 port map( D => 
                           n1446, CK => clk, RN => n306, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_7);
   input_p2_times_b2_div_componentxoutput_sign_gated_reg : DFFRHQX1 port map( D
                           => n4296, CK => clk, RN => n313, Q => 
                           input_p2_times_b2_div_componentxoutput_sign_gated);
   input_times_b0_div_componentxUDxquotient_reg_2 : DFFRHQX1 port map( D => 
                           n1265, CK => clk, RN => n304, Q => 
                           input_times_b0_div_componentxunsigned_output_2);
   output_p2_times_a2_div_componentxUDxquotient_reg_2 : DFFRHQX1 port map( D =>
                           n1384, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_2);
   output_p1_times_a1_div_componentxUDxquotient_reg_2 : DFFRHQX1 port map( D =>
                           n1403, CK => clk, RN => n311, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_2);
   input_p1_times_b1_div_componentxUDxquotient_reg_2 : DFFRHQX1 port map( D => 
                           n1441, CK => clk, RN => n306, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_2);
   input_times_b0_div_componentxUDxquotient_reg_4 : DFFRHQX1 port map( D => 
                           n1267, CK => clk, RN => n304, Q => 
                           input_times_b0_div_componentxunsigned_output_4);
   output_p2_times_a2_div_componentxUDxquotient_reg_4 : DFFRHQX1 port map( D =>
                           n1386, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_4);
   output_p1_times_a1_div_componentxUDxquotient_reg_4 : DFFRHQX1 port map( D =>
                           n1405, CK => clk, RN => n311, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_4);
   input_p1_times_b1_div_componentxUDxquotient_reg_4 : DFFRHQX1 port map( D => 
                           n1443, CK => clk, RN => n306, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_4);
   input_times_b0_div_componentxUDxquotient_reg_1 : DFFRHQX1 port map( D => 
                           n1264, CK => clk, RN => n304, Q => 
                           input_times_b0_div_componentxunsigned_output_1);
   output_p2_times_a2_div_componentxUDxquotient_reg_1 : DFFRHQX1 port map( D =>
                           n1383, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_1);
   output_p1_times_a1_div_componentxUDxquotient_reg_1 : DFFRHQX1 port map( D =>
                           n1402, CK => clk, RN => n311, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_1);
   input_p2_times_b2_div_componentxUDxquotient_reg_1 : DFFRHQX1 port map( D => 
                           n1421, CK => clk, RN => n309, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_1);
   input_times_b0_div_componentxUDxquotient_reg_3 : DFFRHQX1 port map( D => 
                           n1266, CK => clk, RN => n304, Q => 
                           input_times_b0_div_componentxunsigned_output_3);
   output_p2_times_a2_div_componentxUDxquotient_reg_3 : DFFRHQX1 port map( D =>
                           n1385, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_3);
   output_p1_times_a1_div_componentxUDxquotient_reg_3 : DFFRHQX1 port map( D =>
                           n1404, CK => clk, RN => n311, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_3);
   input_p1_times_b1_div_componentxUDxquotient_reg_3 : DFFRHQX1 port map( D => 
                           n1442, CK => clk, RN => n306, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_3);
   input_p2_times_b2_div_componentxUDxquotient_reg_0 : DFFRHQX1 port map( D => 
                           n1420, CK => clk, RN => n309, Q => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_0_port);
   input_times_b0_div_componentxoutput_sign_gated_reg : DFFRHQX1 port map( D =>
                           input_times_b0_div_componentxn62, CK => clk, RN => 
                           n305, Q => 
                           input_times_b0_div_componentxoutput_sign_gated);
   output_p2_times_a2_div_componentxoutput_sign_gated_reg : DFFRHQX1 port map( 
                           D => n4406, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxoutput_sign_gated);
   output_p1_times_a1_div_componentxoutput_sign_gated_reg : DFFRHQX1 port map( 
                           D => n4350, CK => clk, RN => n313, Q => 
                           output_p1_times_a1_div_componentxoutput_sign_gated);
   input_p1_times_b1_div_componentxoutput_sign_gated_reg : DFFRHQX1 port map( D
                           => n4240, CK => clk, RN => n313, Q => 
                           input_p1_times_b1_div_componentxoutput_sign_gated);
   input_p1_times_b1_div_componentxUDxquotient_reg_1 : DFFRHQX1 port map( D => 
                           n1440, CK => clk, RN => n306, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_1);
   input_times_b0_div_componentxUDxquotient_reg_0 : DFFRHQX1 port map( D => 
                           n1263, CK => clk, RN => n304, Q => 
                           input_times_b0_div_componentxunsigned_output_inverted_0_port);
   output_p2_times_a2_div_componentxUDxquotient_reg_0 : DFFRHQX1 port map( D =>
                           n1382, CK => clk, RN => n313, Q => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_0_port);
   output_p1_times_a1_div_componentxUDxquotient_reg_0 : DFFRHQX1 port map( D =>
                           n1401, CK => clk, RN => n311, Q => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_0_port);
   input_p1_times_b1_div_componentxUDxquotient_reg_0 : DFFRHQX1 port map( D => 
                           n1439, CK => clk, RN => n307, Q => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_0_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_0 : 
                           DFFRHQX1 port map( D => change_input_port, CK => clk
                           , RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_0_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_0 : 
                           DFFRHQX1 port map( D => change_input_port, CK => clk
                           , RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_0_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_0 : 
                           DFFRHQX1 port map( D => change_input_port, CK => clk
                           , RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_0_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_0 : 
                           DFFRHQX1 port map( D => change_input_port, CK => clk
                           , RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_0_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_0 : 
                           DFFRHQX1 port map( D => change_input_port, CK => clk
                           , RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_0_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_18 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_17_port, 
                           CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_18_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_17 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_16_port, 
                           CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_17_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_16 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_15_port, 
                           CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_16_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_15 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_14_port, 
                           CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_15_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_14 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_13_port, 
                           CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_14_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_13 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_12_port, 
                           CK => clk, RN => n303, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_13_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_12 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_11_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_12_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_11 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_10_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_11_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_10 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_9_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_10_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_9 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_8_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_9_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_8 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_7_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_8_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_7 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_6_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_7_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_6 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_5_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_6_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_5 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_4_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_5_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_4 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_3_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_4_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_3 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_2_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_3_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_2 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_1_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_2_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_1 : 
                           DFFRHQX1 port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_0_port, 
                           CK => clk, RN => n302, Q => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_1_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_18 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_17_port, 
                           CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_18_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_17 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_16_port, 
                           CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_17_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_16 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_15_port, 
                           CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_16_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_15 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_14_port, 
                           CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_15_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_14 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_13_port, 
                           CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_14_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_13 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_12_port, 
                           CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_13_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_12 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_11_port, 
                           CK => clk, RN => n312, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_12_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_11 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_10_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_11_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_10 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_9_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_10_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_9 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_8_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_9_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_8 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_7_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_8_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_7 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_6_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_7_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_6 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_5_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_6_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_5 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_4_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_5_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_4 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_3_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_4_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_3 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_2_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_3_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_2 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_1_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_2_port);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_1 : 
                           DFFRHQX1 port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_0_port, 
                           CK => clk, RN => n311, Q => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_1_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_18 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_17_port, 
                           CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_18_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_17 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_16_port, 
                           CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_17_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_16 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_15_port, 
                           CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_16_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_15 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_14_port, 
                           CK => clk, RN => n310, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_15_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_14 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_13_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_14_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_13 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_12_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_13_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_12 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_11_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_12_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_11 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_10_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_11_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_10 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_9_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_10_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_9 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_8_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_9_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_8 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_7_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_8_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_7 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_6_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_7_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_6 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_5_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_6_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_5 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_4_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_5_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_4 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_3_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_4_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_3 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_2_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_3_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_2 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_1_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_2_port);
   output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_reg_1 : 
                           DFFRHQX1 port map( D => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_0_port, 
                           CK => clk, RN => n309, Q => 
                           output_p1_times_a1_div_componentxUDxreadiness_propagation_vector_1_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_18 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_17_port, 
                           CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_18_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_17 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_16_port, 
                           CK => clk, RN => n308, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_17_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_16 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_15_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_16_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_15 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_14_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_15_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_14 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_13_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_14_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_13 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_12_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_13_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_12 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_11_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_12_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_11 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_10_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_11_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_10 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_9_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_10_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_9 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_8_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_9_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_8 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_7_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_8_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_7 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_6_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_7_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_6 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_5_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_6_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_5 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_4_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_5_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_4 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_3_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_4_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_3 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_2_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_3_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_2 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_1_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_2_port);
   input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_reg_1 : 
                           DFFRHQX1 port map( D => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_0_port, 
                           CK => clk, RN => n307, Q => 
                           input_p2_times_b2_div_componentxUDxreadiness_propagation_vector_1_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_18 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_17_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_18_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_17 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_16_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_17_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_16 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_15_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_16_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_15 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_14_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_15_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_14 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_13_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_14_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_13 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_12_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_13_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_12 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_11_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_12_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_11 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_10_port, 
                           CK => clk, RN => n290, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_11_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_10 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_9_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_10_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_9 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_8_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_9_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_8 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_7_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_8_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_7 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_6_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_7_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_6 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_5_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_6_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_5 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_4_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_5_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_4 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_3_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_4_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_3 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_2_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_3_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_2 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_1_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_2_port);
   input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_reg_1 : 
                           DFFRHQX1 port map( D => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_0_port, 
                           CK => clk, RN => n289, Q => 
                           input_p1_times_b1_div_componentxUDxreadiness_propagation_vector_1_port);
   input_times_b0_div_componentxUDxreadiness_propagation_vector_reg_19 : DFFRXL
                           port map( D => 
                           input_times_b0_div_componentxUDxreadiness_propagation_vector_18_port, 
                           CK => clk, RN => n283, Q => n8, QN => n257);
   output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_reg_19 : 
                           DFFRXL port map( D => 
                           output_p2_times_a2_div_componentxUDxreadiness_propagation_vector_18_port, 
                           CK => clk, RN => n284, Q => n7, QN => n164);
   U3 : AND2X2 port map( A => change_input_port, B => en, Y => n1);
   U4 : NOR2X1 port map( A => n367, B => n837, Y => n2);
   U5 : NOR2X1 port map( A => n368, B => n996, Y => n3);
   U6 : NOR2X1 port map( A => n367, B => n1155, Y => n4);
   U7 : NOR2X1 port map( A => n368, B => n519, Y => n5);
   U8 : NOR2X1 port map( A => n367, B => n678, Y => n6);
   U9 : NAND2X1 port map( A => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_17_port, B 
                           => n165, Y => n9);
   U10 : NAND2X1 port map( A => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_17_port, B 
                           => input_previous_1_17_port, Y => n10);
   U11 : NAND2X1 port map( A => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_17_port, B 
                           => input_previous_2_17_port, Y => n11);
   U12 : NAND2X1 port map( A => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_17_port, B 
                           => output_previous_2_17_port, Y => n12);
   U13 : NAND2X1 port map( A => 
                           input_times_b0_mul_componentxinput_A_inverted_17_port, B 
                           => input_previous_0_17_port, Y => n13);
   U14 : AND2X2 port map( A => n837, B => en, Y => n14);
   U15 : AND2X2 port map( A => n996, B => en, Y => n15);
   U16 : AND2X2 port map( A => n1155, B => en, Y => n16);
   U17 : AND2X2 port map( A => n519, B => en, Y => n17);
   U18 : AND2X2 port map( A => n678, B => en, Y => n18);
   U19 : AND2X4 port map( A => n25, B => n26, Y => temporary_overflow);
   U20 : NAND2X1 port map( A => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_17_port, B 
                           => n363, Y => n20);
   U21 : NAND2X1 port map( A => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_17_port, B 
                           => n336, Y => n21);
   U22 : NAND2X1 port map( A => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_17_port, B 
                           => n327, Y => n22);
   U23 : NAND2X1 port map( A => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_17_port, B 
                           => n354, Y => n23);
   U24 : NAND2X1 port map( A => 
                           input_times_b0_mul_componentxinput_B_inverted_17_port, B 
                           => n345, Y => n24);
   U25 : NAND2X1 port map( A => output_contracterxn1, B => output_contracterxn2
                           , Y => n25);
   U26 : NAND2X1 port map( A => n27, B => n28, Y => n26);
   U27 : INVX1 port map( A => output_contracterxn4, Y => n27);
   U28 : INVX1 port map( A => output_contracterxn3, Y => n28);
   U29 : XNOR2X4 port map( A => n79, B => n4168, Y => output_signal_1_port);
   U30 : INVXL port map( A => output_signal_1_port, Y => n1226);
   U31 : INVX1 port map( A => n348, Y => n343);
   U32 : INVX1 port map( A => n342, Y => n340);
   U33 : INVX1 port map( A => n333, Y => n331);
   U34 : INVX1 port map( A => n324, Y => n322);
   U35 : INVX1 port map( A => n360, Y => n358);
   U36 : INVX1 port map( A => n351, Y => n349);
   U37 : INVX1 port map( A => en, Y => n370);
   U38 : INVX1 port map( A => en, Y => n369);
   U39 : INVX1 port map( A => en, Y => n372);
   U40 : INVX1 port map( A => en, Y => n371);
   U41 : INVX1 port map( A => en, Y => n367);
   U42 : NOR2BX1 port map( AN => n3817, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_15,
                           Y => n3816);
   U43 : NAND2BX1 port map( AN => 
                           output_p1_times_a1_mul_componentxunsigned_output_16,
                           B => n3816, Y => n3815);
   U44 : INVX1 port map( A => 
                           output_p1_times_a1_mul_componentxunsigned_output_9, 
                           Y => n462);
   U45 : NOR2BX1 port map( AN => n3721, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_15, 
                           Y => n3720);
   U46 : NOR2BX1 port map( AN => n3673, B => 
                           input_times_b0_mul_componentxunsigned_output_15, Y 
                           => n3672);
   U47 : NAND2BX1 port map( AN => 
                           input_p1_times_b1_mul_componentxunsigned_output_16, 
                           B => n3720, Y => n3719);
   U48 : NAND2BX1 port map( AN => 
                           input_p2_times_b2_mul_componentxunsigned_output_16, 
                           B => n3768, Y => n3767);
   U49 : NAND2BX1 port map( AN => 
                           output_p2_times_a2_mul_componentxunsigned_output_16,
                           B => n3864, Y => n3863);
   U50 : NAND2BX1 port map( AN => 
                           input_times_b0_mul_componentxunsigned_output_16, B 
                           => n3672, Y => n3671);
   U51 : NOR2BX1 port map( AN => n3769, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_15, 
                           Y => n3768);
   U52 : NOR2BX1 port map( AN => n3865, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_15,
                           Y => n3864);
   U53 : INVX1 port map( A => input_p1_times_b1_mul_componentxunsigned_output_9
                           , Y => n939);
   U54 : INVX1 port map( A => input_p2_times_b2_mul_componentxunsigned_output_9
                           , Y => n1098);
   U55 : INVX1 port map( A => 
                           output_p2_times_a2_mul_componentxunsigned_output_9, 
                           Y => n621);
   U56 : INVX1 port map( A => input_times_b0_mul_componentxunsigned_output_9, Y
                           => n780);
   U57 : NOR3X1 port map( A => 
                           output_p1_times_a1_mul_componentxunsigned_output_13,
                           B => 
                           output_p1_times_a1_mul_componentxunsigned_output_14,
                           C => n3818, Y => n3817);
   U58 : XOR2X1 port map( A => n2360, B => n2361, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_14)
                           ;
   U59 : XOR2X1 port map( A => n2356, B => n2357, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_16)
                           ;
   U60 : XOR2X1 port map( A => n2362, B => n2363, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_13)
                           ;
   U61 : XOR2X1 port map( A => n2349, B => n2350, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_9);
   U62 : XOR2X1 port map( A => n2366, B => n2367, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_11)
                           ;
   U63 : XOR2X1 port map( A => n2358, B => n2359, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_15)
                           ;
   U64 : XOR2X1 port map( A => n2351, B => n2352, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_8);
   U65 : XOR2X1 port map( A => n2364, B => n2365, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_12)
                           ;
   U66 : XOR2X1 port map( A => n2368, B => n2369, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_10)
                           ;
   U67 : XOR2X1 port map( A => n2316, B => n2317, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_15);
   U68 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn518
                           , B => 
                           input_times_b0_mul_componentxUMxAdder_finalxn519, Y 
                           => input_times_b0_mul_componentxunsigned_output_15);
   U69 : XOR2X1 port map( A => n2314, B => n2315, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_16);
   U70 : XOR2X1 port map( A => n2335, B => n2336, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_16);
   U71 : XOR2X1 port map( A => n2377, B => n2378, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_16)
                           ;
   U72 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn496
                           , B => 
                           input_times_b0_mul_componentxUMxAdder_finalxn497, Y 
                           => input_times_b0_mul_componentxunsigned_output_16);
   U73 : NOR3X1 port map( A => 
                           input_p1_times_b1_mul_componentxunsigned_output_13, 
                           B => 
                           input_p1_times_b1_mul_componentxunsigned_output_14, 
                           C => n3722, Y => n3721);
   U74 : NOR3X1 port map( A => 
                           input_p2_times_b2_mul_componentxunsigned_output_13, 
                           B => 
                           input_p2_times_b2_mul_componentxunsigned_output_14, 
                           C => n3770, Y => n3769);
   U75 : NOR3X1 port map( A => 
                           output_p2_times_a2_mul_componentxunsigned_output_13,
                           B => 
                           output_p2_times_a2_mul_componentxunsigned_output_14,
                           C => n3866, Y => n3865);
   U76 : NOR3X1 port map( A => input_times_b0_mul_componentxunsigned_output_13,
                           B => input_times_b0_mul_componentxunsigned_output_14
                           , C => n3674, Y => n3673);
   U77 : XOR2X1 port map( A => n2320, B => n2321, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_13);
   U78 : XOR2X1 port map( A => n2341, B => n2342, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_13);
   U79 : XOR2X1 port map( A => n2383, B => n2384, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_13)
                           ;
   U80 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn562
                           , B => 
                           input_times_b0_mul_componentxUMxAdder_finalxn563, Y 
                           => input_times_b0_mul_componentxunsigned_output_13);
   U81 : XOR2X1 port map( A => n2307, B => n2308, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_9);
   U82 : XOR2X1 port map( A => n2328, B => n2329, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_9);
   U83 : XOR2X1 port map( A => n2370, B => n2371, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_9);
   U84 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn2, 
                           B => input_times_b0_mul_componentxUMxAdder_finalxn3,
                           Y => input_times_b0_mul_componentxunsigned_output_9)
                           ;
   U85 : XOR2X1 port map( A => n2324, B => n2325, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_11);
   U86 : XOR2X1 port map( A => n2345, B => n2346, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_11);
   U87 : XOR2X1 port map( A => n2387, B => n2388, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_11)
                           ;
   U88 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn606
                           , B => 
                           input_times_b0_mul_componentxUMxAdder_finalxn607, Y 
                           => input_times_b0_mul_componentxunsigned_output_11);
   U89 : XOR2X1 port map( A => n2337, B => n2338, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_15);
   U90 : XOR2X1 port map( A => n2379, B => n2380, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_15)
                           ;
   U91 : XOR2X1 port map( A => n2309, B => n2310, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_8);
   U92 : XOR2X1 port map( A => n2318, B => n2319, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_14);
   U93 : XOR2X1 port map( A => n2330, B => n2331, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_8);
   U94 : XOR2X1 port map( A => n2339, B => n2340, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_14);
   U95 : XOR2X1 port map( A => n2372, B => n2373, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_8);
   U96 : XOR2X1 port map( A => n2381, B => n2382, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_14)
                           ;
   U97 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn24,
                           B => input_times_b0_mul_componentxUMxAdder_finalxn25
                           , Y => 
                           input_times_b0_mul_componentxunsigned_output_8);
   U98 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn540
                           , B => 
                           input_times_b0_mul_componentxUMxAdder_finalxn541, Y 
                           => input_times_b0_mul_componentxunsigned_output_14);
   U99 : XOR2X1 port map( A => n2322, B => n2323, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_12);
   U100 : XOR2X1 port map( A => n2343, B => n2344, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_12);
   U101 : XOR2X1 port map( A => n2385, B => n2386, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_12)
                           ;
   U102 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxAdder_finalxn584, B 
                           => input_times_b0_mul_componentxUMxAdder_finalxn585,
                           Y => input_times_b0_mul_componentxunsigned_output_12
                           );
   U103 : XOR2X1 port map( A => n2326, B => n2327, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_10);
   U104 : XOR2X1 port map( A => n2347, B => n2348, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_10);
   U105 : XOR2X1 port map( A => n2389, B => n2390, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_10)
                           ;
   U106 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxAdder_finalxn628, B 
                           => input_times_b0_mul_componentxUMxAdder_finalxn629,
                           Y => input_times_b0_mul_componentxunsigned_output_10
                           );
   U107 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_9_port, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_9_port, 
                           B0 => n2349, B1 => n2350, Y => n2369);
   U108 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_11_port, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_11_port, 
                           B0 => n2366, B1 => n2367, Y => n2365);
   U109 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_13_port, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_13_port, 
                           B0 => n2362, B1 => n2363, Y => n2361);
   U110 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_15_port, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_15_port, 
                           B0 => n2358, B1 => n2359, Y => n2357);
   U111 : OAI2BB2X1 port map( B0 => n2365, B1 => n2364, A0N => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_12_port, 
                           A1N => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_12_port, Y 
                           => n2362);
   U112 : OAI2BB2X1 port map( B0 => n2361, B1 => n2360, A0N => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_14_port, 
                           A1N => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_14_port, Y 
                           => n2358);
   U113 : OAI2BB2X1 port map( B0 => n2369, B1 => n2368, A0N => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_10_port, 
                           A1N => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_10_port, Y 
                           => n2366);
   U114 : OAI2BB2X1 port map( B0 => n2352, B1 => n2351, A0N => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_8_port, 
                           A1N => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_8_port, Y 
                           => n2349);
   U115 : OAI2BB2X1 port map( B0 => n2357, B1 => n2356, A0N => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_16_port, 
                           A1N => n407, Y => n2354);
   U116 : XNOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_8_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_8_port, Y 
                           => n2351);
   U117 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_7_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_7_port, Y 
                           => n2353);
   U118 : NAND2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_7_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_7_port, Y 
                           => n2352);
   U119 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128220800_128221024_128221136, B 
                           => n3320, Y => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_15_port);
   U120 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_9_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_9_port, Y 
                           => n2350);
   U121 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_11_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_11_port, Y 
                           => n2367);
   U122 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_13_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_13_port, Y 
                           => n2363);
   U123 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_15_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_15_port, Y 
                           => n2359);
   U124 : OR3XL port map( A => 
                           output_p1_times_a1_mul_componentxunsigned_output_11,
                           B => 
                           output_p1_times_a1_mul_componentxunsigned_output_12,
                           C => n3820, Y => n3818);
   U125 : XNOR2X1 port map( A => n407, B => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_16_port, Y 
                           => n2356);
   U126 : XNOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_10_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_10_port, Y 
                           => n2368);
   U127 : XNOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_12_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_12_port, Y 
                           => n2364);
   U128 : XNOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_14_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_14_port, Y 
                           => n2360);
   U129 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128315464_128315632_128315800, B 
                           => n3322, Y => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_16_port);
   U130 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_13_port, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_13_port, 
                           B0 => n2320, B1 => n2321, Y => n2319);
   U131 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsecond_vector_13_port, 
                           A1 => 
                           input_times_b0_mul_componentxUMxfirst_vector_13_port
                           , B0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn562, B1
                           => input_times_b0_mul_componentxUMxAdder_finalxn563,
                           Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn541);
   U132 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_15_port, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_15_port, 
                           B0 => n2316, B1 => n2317, Y => n2315);
   U133 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_15_port, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_15_port, 
                           B0 => n2337, B1 => n2338, Y => n2336);
   U134 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_15_port, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_15_port, 
                           B0 => n2379, B1 => n2380, Y => n2378);
   U135 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsecond_vector_15_port, 
                           A1 => 
                           input_times_b0_mul_componentxUMxfirst_vector_15_port
                           , B0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn518, B1
                           => input_times_b0_mul_componentxUMxAdder_finalxn519,
                           Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn497);
   U136 : OAI2BB2X1 port map( B0 => n2319, B1 => n2318, A0N => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_14_port, 
                           A1N => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_14_port, Y 
                           => n2316);
   U137 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn541, B1
                           => input_times_b0_mul_componentxUMxAdder_finalxn540,
                           A0N => 
                           input_times_b0_mul_componentxUMxsecond_vector_14_port, 
                           A1N => 
                           input_times_b0_mul_componentxUMxfirst_vector_14_port
                           , Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn518);
   U138 : OAI2BB2X1 port map( B0 => n2315, B1 => n2314, A0N => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_16_port, 
                           A1N => n883, Y => n2312);
   U139 : OAI2BB2X1 port map( B0 => n2336, B1 => n2335, A0N => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_16_port, 
                           A1N => n1042, Y => n2333);
   U140 : OAI2BB2X1 port map( B0 => n2378, B1 => n2377, A0N => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_16_port, 
                           A1N => n565, Y => n2375);
   U141 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn497, B1
                           => input_times_b0_mul_componentxUMxAdder_finalxn496,
                           A0N => 
                           input_times_b0_mul_componentxUMxsecond_vector_16_port, 
                           A1N => n724, Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn474);
   U142 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128220800_128221024_128221136, B 
                           => n2852, Y => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_15_port);
   U143 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128220800_128221024_128221136, B 
                           => n3086, Y => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_15_port);
   U144 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128220800_128221024_128221136, B 
                           => n3554, Y => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_15_port);
   U145 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128220800_128221024_128221136, B 
                           => n2618, Y => 
                           input_times_b0_mul_componentxUMxsecond_vector_15_port);
   U146 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_13_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_13_port, Y 
                           => n2321);
   U147 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_13_port
                           , B => 
                           input_times_b0_mul_componentxUMxsecond_vector_13_port, Y 
                           => input_times_b0_mul_componentxUMxAdder_finalxn563)
                           ;
   U148 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_15_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_15_port, Y 
                           => n2317);
   U149 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_15_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_15_port, Y 
                           => n2338);
   U150 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_15_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_15_port, Y 
                           => n2380);
   U151 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_15_port
                           , B => 
                           input_times_b0_mul_componentxUMxsecond_vector_15_port, Y 
                           => input_times_b0_mul_componentxUMxAdder_finalxn519)
                           ;
   U152 : XNOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_14_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_14_port, Y 
                           => n2318);
   U153 : XNOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_14_port
                           , B => 
                           input_times_b0_mul_componentxUMxsecond_vector_14_port, Y 
                           => input_times_b0_mul_componentxUMxAdder_finalxn540)
                           ;
   U154 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_9_port, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_9_port, 
                           B0 => n2307, B1 => n2308, Y => n2327);
   U155 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_9_port, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_9_port, 
                           B0 => n2328, B1 => n2329, Y => n2348);
   U156 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_9_port, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_9_port, 
                           B0 => n2370, B1 => n2371, Y => n2390);
   U157 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsecond_vector_9_port
                           , A1 => 
                           input_times_b0_mul_componentxUMxfirst_vector_9_port,
                           B0 => input_times_b0_mul_componentxUMxAdder_finalxn2
                           , B1 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn3, Y =>
                           input_times_b0_mul_componentxUMxAdder_finalxn629);
   U158 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_11_port, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_11_port, 
                           B0 => n2324, B1 => n2325, Y => n2323);
   U159 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_11_port, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_11_port, 
                           B0 => n2345, B1 => n2346, Y => n2344);
   U160 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_11_port, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_11_port, 
                           B0 => n2387, B1 => n2388, Y => n2386);
   U161 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsecond_vector_11_port, 
                           A1 => 
                           input_times_b0_mul_componentxUMxfirst_vector_11_port
                           , B0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn606, B1
                           => input_times_b0_mul_componentxUMxAdder_finalxn607,
                           Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn585);
   U162 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_13_port, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_13_port, 
                           B0 => n2341, B1 => n2342, Y => n2340);
   U163 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_13_port, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_13_port, 
                           B0 => n2383, B1 => n2384, Y => n2382);
   U164 : OAI2BB2X1 port map( B0 => n2323, B1 => n2322, A0N => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_12_port, 
                           A1N => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_12_port, Y 
                           => n2320);
   U165 : OAI2BB2X1 port map( B0 => n2344, B1 => n2343, A0N => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_12_port, 
                           A1N => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_12_port, Y 
                           => n2341);
   U166 : OAI2BB2X1 port map( B0 => n2386, B1 => n2385, A0N => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_12_port, 
                           A1N => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_12_port, Y 
                           => n2383);
   U167 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn585, B1
                           => input_times_b0_mul_componentxUMxAdder_finalxn584,
                           A0N => 
                           input_times_b0_mul_componentxUMxsecond_vector_12_port, 
                           A1N => 
                           input_times_b0_mul_componentxUMxfirst_vector_12_port
                           , Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn562);
   U168 : OAI2BB2X1 port map( B0 => n2340, B1 => n2339, A0N => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_14_port, 
                           A1N => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_14_port, Y 
                           => n2337);
   U169 : OAI2BB2X1 port map( B0 => n2382, B1 => n2381, A0N => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_14_port, 
                           A1N => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_14_port, Y 
                           => n2379);
   U170 : OAI2BB2X1 port map( B0 => n2327, B1 => n2326, A0N => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_10_port, 
                           A1N => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_10_port, Y 
                           => n2324);
   U171 : OAI2BB2X1 port map( B0 => n2348, B1 => n2347, A0N => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_10_port, 
                           A1N => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_10_port, Y 
                           => n2345);
   U172 : OAI2BB2X1 port map( B0 => n2390, B1 => n2389, A0N => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_10_port, 
                           A1N => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_10_port, Y 
                           => n2387);
   U173 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn629, B1
                           => input_times_b0_mul_componentxUMxAdder_finalxn628,
                           A0N => 
                           input_times_b0_mul_componentxUMxsecond_vector_10_port, 
                           A1N => 
                           input_times_b0_mul_componentxUMxfirst_vector_10_port
                           , Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn606);
   U174 : OAI2BB2X1 port map( B0 => n2310, B1 => n2309, A0N => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_8_port, 
                           A1N => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_8_port, Y 
                           => n2307);
   U175 : OAI2BB2X1 port map( B0 => n2331, B1 => n2330, A0N => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_8_port, 
                           A1N => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_8_port, Y 
                           => n2328);
   U176 : OAI2BB2X1 port map( B0 => n2373, B1 => n2372, A0N => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_8_port, 
                           A1N => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_8_port, Y 
                           => n2370);
   U177 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn25, B1 
                           => input_times_b0_mul_componentxUMxAdder_finalxn24, 
                           A0N => 
                           input_times_b0_mul_componentxUMxsecond_vector_8_port
                           , A1N => 
                           input_times_b0_mul_componentxUMxfirst_vector_8_port,
                           Y => input_times_b0_mul_componentxUMxAdder_finalxn2)
                           ;
   U178 : NAND2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_7_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_7_port, Y 
                           => n2310);
   U179 : NAND2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_7_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_7_port, Y 
                           => n2331);
   U180 : NAND2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_7_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_7_port, Y 
                           => n2373);
   U181 : NAND2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsecond_vector_7_port
                           , B => 
                           input_times_b0_mul_componentxUMxfirst_vector_7_port,
                           Y => input_times_b0_mul_componentxUMxAdder_finalxn25
                           );
   U182 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_9_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_9_port, Y 
                           => n2308);
   U183 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_9_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_9_port, Y 
                           => n2329);
   U184 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_9_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_9_port, Y 
                           => n2371);
   U185 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_9_port,
                           B => 
                           input_times_b0_mul_componentxUMxsecond_vector_9_port
                           , Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn3);
   U186 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_11_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_11_port, Y 
                           => n2325);
   U187 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_11_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_11_port, Y 
                           => n2346);
   U188 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_11_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_11_port, Y 
                           => n2388);
   U189 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_11_port
                           , B => 
                           input_times_b0_mul_componentxUMxsecond_vector_11_port, Y 
                           => input_times_b0_mul_componentxUMxAdder_finalxn607)
                           ;
   U190 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_13_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_13_port, Y 
                           => n2342);
   U191 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_13_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_13_port, Y 
                           => n2384);
   U192 : OR3XL port map( A => 
                           input_p1_times_b1_mul_componentxunsigned_output_11, 
                           B => 
                           input_p1_times_b1_mul_componentxunsigned_output_12, 
                           C => n3724, Y => n3722);
   U193 : OR3XL port map( A => 
                           input_p2_times_b2_mul_componentxunsigned_output_11, 
                           B => 
                           input_p2_times_b2_mul_componentxunsigned_output_12, 
                           C => n3772, Y => n3770);
   U194 : OR3XL port map( A => 
                           output_p2_times_a2_mul_componentxunsigned_output_11,
                           B => 
                           output_p2_times_a2_mul_componentxunsigned_output_12,
                           C => n3868, Y => n3866);
   U195 : OR3XL port map( A => input_times_b0_mul_componentxunsigned_output_11,
                           B => input_times_b0_mul_componentxunsigned_output_12
                           , C => n3676, Y => n3674);
   U196 : XNOR2X1 port map( A => n883, B => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_16_port, Y 
                           => n2314);
   U197 : XNOR2X1 port map( A => n1042, B => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_16_port, Y 
                           => n2335);
   U198 : XNOR2X1 port map( A => n565, B => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_16_port, Y 
                           => n2377);
   U199 : XNOR2X1 port map( A => n724, B => 
                           input_times_b0_mul_componentxUMxsecond_vector_16_port, Y 
                           => input_times_b0_mul_componentxUMxAdder_finalxn496)
                           ;
   U200 : XNOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_8_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_8_port, Y 
                           => n2309);
   U201 : XNOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_8_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_8_port, Y 
                           => n2330);
   U202 : XNOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_8_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_8_port, Y 
                           => n2372);
   U203 : XNOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_8_port,
                           B => 
                           input_times_b0_mul_componentxUMxsecond_vector_8_port
                           , Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn24);
   U204 : XNOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_10_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_10_port, Y 
                           => n2326);
   U205 : XNOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_10_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_10_port, Y 
                           => n2347);
   U206 : XNOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_10_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_10_port, Y 
                           => n2389);
   U207 : XNOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_10_port
                           , B => 
                           input_times_b0_mul_componentxUMxsecond_vector_10_port, Y 
                           => input_times_b0_mul_componentxUMxAdder_finalxn628)
                           ;
   U208 : XNOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_12_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_12_port, Y 
                           => n2322);
   U209 : XNOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_12_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_12_port, Y 
                           => n2343);
   U210 : XNOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_12_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_12_port, Y 
                           => n2385);
   U211 : XNOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_12_port
                           , B => 
                           input_times_b0_mul_componentxUMxsecond_vector_12_port, Y 
                           => input_times_b0_mul_componentxUMxAdder_finalxn584)
                           ;
   U212 : XNOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_14_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_14_port, Y 
                           => n2339);
   U213 : XNOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_14_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_14_port, Y 
                           => n2381);
   U214 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128315464_128315632_128315800, B 
                           => n2854, Y => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_16_port);
   U215 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128315464_128315632_128315800, B 
                           => n3088, Y => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_16_port);
   U216 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128315464_128315632_128315800, B 
                           => n3556, Y => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_16_port);
   U217 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128315464_128315632_128315800, B 
                           => n2620, Y => 
                           input_times_b0_mul_componentxUMxsecond_vector_16_port);
   U218 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_7_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_7_port, Y 
                           => n2311);
   U219 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_7_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_7_port, Y 
                           => n2332);
   U220 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_7_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_7_port, Y 
                           => n2374);
   U221 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_7_port,
                           B => 
                           input_times_b0_mul_componentxUMxsecond_vector_7_port
                           , Y => 
                           input_times_b0_mul_componentxUMxAdder_finalxn47);
   U222 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_8_port);
   U223 : NAND3BX1 port map( AN => 
                           output_p1_times_a1_mul_componentxunsigned_output_10,
                           B => n462, C => n3807, Y => n3820);
   U224 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_6_port);
   U225 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_9_port);
   U226 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n452, Y => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_11_port);
   U227 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n431, Y => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_13_port);
   U228 : XOR2X1 port map( A => n429, B => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128262496_128126088_128126312, Y 
                           => n3313);
   U229 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126816_128126928, B 
                           => n416, Y => n3320);
   U230 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128237920_128238088, B 
                           => n414, Y => n3322);
   U231 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_7_port);
   U232 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_10_port);
   U233 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n440, Y => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_12_port);
   U234 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n422, Y => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_14_port);
   U235 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128263168_128126424_128126648, B 
                           => n3315, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128220800_128221024_128221136);
   U236 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_9_port);
   U237 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_11_port);
   U238 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n440, Y => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_13_port);
   U239 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_7_port);
   U240 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124744_128124968_128125136, B 
                           => n3305, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125248_128219960_128220240);
   U241 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125080_128125304_128125472, B 
                           => n3307, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125584_128220184_128220408);
   U242 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125416_128125640_128125808, B 
                           => n3309, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125920_128220352_128220576);
   U243 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125752_128125976_128126144, B 
                           => n3311, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128126256_128220520_128220744);
   U244 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126480_128126592, B 
                           => n3313, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128220688_128220856_128220968);
   U245 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_8_port);
   U246 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_10_port);
   U247 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n452, Y => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_12_port);
   U248 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n431, Y => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_14_port);
   U249 : INVX1 port map( A => n3314, Y => n416);
   U250 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
                           A1 => n429, B0 => n3313, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126480_128126592, Y 
                           => n3314);
   U251 : INVX1 port map( A => n3321, Y => n407);
   U252 : AOI22X1 port map( A0 => n416, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126816_128126928, 
                           B0 => n3320, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128220800_128221024_128221136, Y 
                           => n3321);
   U253 : AOI22X1 port map( A0 => n414, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128237920_128238088, 
                           B0 => n3322, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128315464_128315632_128315800, Y 
                           => n3323);
   U254 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126760_128237640_128237808, B 
                           => n3317, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128315464_128315632_128315800);
   U255 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n422, Y => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_15_port);
   U256 : INVX1 port map( A => n2846, Y => n892);
   U257 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
                           A1 => n905, B0 => n2845, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126480_128126592, Y 
                           => n2846);
   U258 : INVX1 port map( A => n2612, Y => n733);
   U259 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
                           A1 => n746, B0 => n2611, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126480_128126592, Y 
                           => n2612);
   U260 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n907, Y => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_13_port);
   U261 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n748, Y => 
                           input_times_b0_mul_componentxUMxsecond_vector_13_port);
   U262 : XOR2X1 port map( A => n905, B => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128262496_128126088_128126312, Y 
                           => n2845);
   U263 : XOR2X1 port map( A => n1064, B => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128262496_128126088_128126312, Y 
                           => n3079);
   U264 : XOR2X1 port map( A => n587, B => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128262496_128126088_128126312, Y 
                           => n3547);
   U265 : XOR2X1 port map( A => n746, B => 
                           input_times_b0_mul_componentxUMxsum_layer4_128262496_128126088_128126312, Y 
                           => n2611);
   U266 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126816_128126928, B 
                           => n892, Y => n2852);
   U267 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126816_128126928, B 
                           => n1051, Y => n3086);
   U268 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126816_128126928, B 
                           => n574, Y => n3554);
   U269 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126816_128126928, B 
                           => n733, Y => n2618);
   U270 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n898, Y => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_14_port);
   U271 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n739, Y => 
                           input_times_b0_mul_componentxUMxsecond_vector_14_port);
   U272 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125752_128125976_128126144, B 
                           => n2843, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128126256_128220520_128220744);
   U273 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125752_128125976_128126144, B 
                           => n2609, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128126256_128220520_128220744);
   U274 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126480_128126592, B 
                           => n2845, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128220688_128220856_128220968);
   U275 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126480_128126592, B 
                           => n2611, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128220688_128220856_128220968);
   U276 : INVX1 port map( A => n3080, Y => n1051);
   U277 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
                           A1 => n1064, B0 => n3079, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126480_128126592, Y 
                           => n3080);
   U278 : INVX1 port map( A => n3548, Y => n574);
   U279 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128262496_128126088_128126312, 
                           A1 => n587, B0 => n3547, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126480_128126592, Y 
                           => n3548);
   U280 : AOI22X1 port map( A0 => n890, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128237920_128238088, 
                           B0 => n2854, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128315464_128315632_128315800, Y 
                           => n2855);
   U281 : AOI22X1 port map( A0 => n1049, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128237920_128238088, 
                           B0 => n3088, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128315464_128315632_128315800, Y 
                           => n3089);
   U282 : AOI22X1 port map( A0 => n572, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128237920_128238088, 
                           B0 => n3556, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128315464_128315632_128315800, Y 
                           => n3557);
   U283 : AOI22X1 port map( A0 => n731, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128237920_128238088, 
                           B0 => n2620, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer5_128315464_128315632_128315800, Y 
                           => n2621);
   U284 : NAND3BX1 port map( AN => 
                           input_p1_times_b1_mul_componentxunsigned_output_10, 
                           B => n939, C => n3711, Y => n3724);
   U285 : NAND3BX1 port map( AN => 
                           input_p2_times_b2_mul_componentxunsigned_output_10, 
                           B => n1098, C => n3759, Y => n3772);
   U286 : NAND3BX1 port map( AN => 
                           output_p2_times_a2_mul_componentxunsigned_output_10,
                           B => n621, C => n3855, Y => n3868);
   U287 : NAND3BX1 port map( AN => 
                           input_times_b0_mul_componentxunsigned_output_10, B 
                           => n780, C => n3663, Y => n3676);
   U288 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_9_port);
   U289 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_9_port);
   U290 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_9_port);
   U291 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           input_times_b0_mul_componentxUMxsecond_vector_9_port
                           );
   U292 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n929, Y => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_11_port);
   U293 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n1088, Y => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_11_port);
   U294 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n611, Y => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_11_port);
   U295 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n770, Y => 
                           input_times_b0_mul_componentxUMxsecond_vector_11_port);
   U296 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n1066, Y => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_13_port);
   U297 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n589, Y => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_13_port);
   U298 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128237920_128238088, B 
                           => n890, Y => n2854);
   U299 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128237920_128238088, B 
                           => n1049, Y => n3088);
   U300 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128237920_128238088, B 
                           => n572, Y => n3556);
   U301 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128237920_128238088, B 
                           => n731, Y => n2620);
   U302 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_7_port);
   U303 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_7_port);
   U304 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_7_port);
   U305 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           input_times_b0_mul_componentxUMxsecond_vector_7_port
                           );
   U306 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_8_port);
   U307 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_8_port);
   U308 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_8_port);
   U309 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           input_times_b0_mul_componentxUMxsecond_vector_8_port
                           );
   U310 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_10_port);
   U311 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_10_port);
   U312 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_10_port);
   U313 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           input_times_b0_mul_componentxUMxsecond_vector_10_port);
   U314 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n916, Y => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_12_port);
   U315 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n1075, Y => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_12_port);
   U316 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n598, Y => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_12_port);
   U317 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n757, Y => 
                           input_times_b0_mul_componentxUMxsecond_vector_12_port);
   U318 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n1057, Y => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_14_port);
   U319 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n580, Y => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_14_port);
   U320 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128263168_128126424_128126648, B 
                           => n2847, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128220800_128221024_128221136);
   U321 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128263168_128126424_128126648, B 
                           => n3081, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128220800_128221024_128221136);
   U322 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128263168_128126424_128126648, B 
                           => n3549, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128220800_128221024_128221136);
   U323 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128263168_128126424_128126648, B 
                           => n2613, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128220800_128221024_128221136);
   U324 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126760_128237640_128237808, B 
                           => n2849, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128315464_128315632_128315800);
   U325 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126760_128237640_128237808, B 
                           => n3083, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128315464_128315632_128315800);
   U326 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126760_128237640_128237808, B 
                           => n3551, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128315464_128315632_128315800);
   U327 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126760_128237640_128237808, B 
                           => n2615, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128315464_128315632_128315800);
   U328 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_9_port);
   U329 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_9_port);
   U330 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_9_port);
   U331 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219624_128219848, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219456_128219680, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_9_port)
                           ;
   U332 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_11_port);
   U333 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_11_port);
   U334 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_11_port);
   U335 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125248_128219960_128220240, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219792_128220016, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_11_port
                           );
   U336 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n916, Y => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_13_port);
   U337 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n1075, Y => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_13_port);
   U338 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n598, Y => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_13_port);
   U339 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125920_128220352_128220576, B 
                           => n757, Y => 
                           input_times_b0_mul_componentxUMxfirst_vector_13_port
                           );
   U340 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n898, Y => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_15_port);
   U341 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n1057, Y => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_15_port);
   U342 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n580, Y => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_15_port);
   U343 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128220688_128220856_128220968, B 
                           => n739, Y => 
                           input_times_b0_mul_componentxUMxfirst_vector_15_port
                           );
   U344 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_7_port);
   U345 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_7_port)
                           ;
   U346 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124744_128124968_128125136, B 
                           => n2837, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125248_128219960_128220240);
   U347 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124744_128124968_128125136, B 
                           => n3071, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125248_128219960_128220240);
   U348 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124744_128124968_128125136, B 
                           => n3539, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125248_128219960_128220240);
   U349 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124744_128124968_128125136, B 
                           => n2603, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125248_128219960_128220240);
   U350 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125080_128125304_128125472, B 
                           => n2839, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125584_128220184_128220408);
   U351 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125080_128125304_128125472, B 
                           => n3073, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125584_128220184_128220408);
   U352 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125080_128125304_128125472, B 
                           => n3541, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125584_128220184_128220408);
   U353 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125080_128125304_128125472, B 
                           => n2605, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125584_128220184_128220408);
   U354 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125416_128125640_128125808, B 
                           => n2841, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125920_128220352_128220576);
   U355 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125416_128125640_128125808, B 
                           => n3075, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125920_128220352_128220576);
   U356 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125416_128125640_128125808, B 
                           => n3543, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125920_128220352_128220576);
   U357 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125416_128125640_128125808, B 
                           => n2607, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125920_128220352_128220576);
   U358 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125752_128125976_128126144, B 
                           => n3077, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128126256_128220520_128220744);
   U359 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125752_128125976_128126144, B 
                           => n3545, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128126256_128220520_128220744);
   U360 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126480_128126592, B 
                           => n3079, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128220688_128220856_128220968);
   U361 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126480_128126592, B 
                           => n3547, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128220688_128220856_128220968);
   U362 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_8_port);
   U363 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_8_port);
   U364 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_8_port);
   U365 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219456_128219680, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219288_128219512, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_8_port)
                           ;
   U366 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_10_port);
   U367 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_10_port);
   U368 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_10_port);
   U369 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219792_128220016, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219624_128219848, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_10_port
                           );
   U370 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n929, Y => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_12_port);
   U371 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n1088, Y => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_12_port);
   U372 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n611, Y => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_12_port);
   U373 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128125584_128220184_128220408, B 
                           => n770, Y => 
                           input_times_b0_mul_componentxUMxfirst_vector_12_port
                           );
   U374 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n907, Y => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_14_port);
   U375 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n1066, Y => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_14_port);
   U376 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n589, Y => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_14_port);
   U377 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128126256_128220520_128220744, B 
                           => n748, Y => 
                           input_times_b0_mul_componentxUMxfirst_vector_14_port
                           );
   U378 : INVX1 port map( A => n2853, Y => n883);
   U379 : AOI22X1 port map( A0 => n892, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126816_128126928, 
                           B0 => n2852, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128220800_128221024_128221136, Y 
                           => n2853);
   U380 : INVX1 port map( A => n3087, Y => n1042);
   U381 : AOI22X1 port map( A0 => n1051, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126816_128126928, 
                           B0 => n3086, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128220800_128221024_128221136, Y 
                           => n3087);
   U382 : INVX1 port map( A => n3555, Y => n565);
   U383 : AOI22X1 port map( A0 => n574, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126816_128126928, 
                           B0 => n3554, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128220800_128221024_128221136, Y 
                           => n3555);
   U384 : INVX1 port map( A => n2619, Y => n724);
   U385 : AOI22X1 port map( A0 => n733, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126816_128126928, 
                           B0 => n2618, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer5_128220800_128221024_128221136, Y 
                           => n2619);
   U386 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_6_port);
   U387 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_6_port);
   U388 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_6_port);
   U389 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_6_port)
                           ;
   U390 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_7_port);
   U391 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219288_128219512, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219120_128219344, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_7_port);
   U392 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219456_128219680);
   U393 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246952_128247176_128247344, B 
                           => n3285, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128247456_128124464_128124688);
   U394 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246616_128246840_128247008, B 
                           => n3283, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128247120_128124240_128124520);
   U395 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n481, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219624_128219848);
   U396 : BUFX3 port map( A => n398, Y => n112);
   U397 : BUFX3 port map( A => n398, Y => n111);
   U398 : NOR3X1 port map( A => output_signal_7_port, B => 
                           output_previous_1_8_port, C => n3777, Y => n3775);
   U399 : NOR3X1 port map( A => n2353, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_8, 
                           C => n3809, Y => n3807);
   U400 : NAND3BX1 port map( AN => output_previous_1_10_port, B => n1210, C => 
                           n3775, Y => n3788);
   U401 : INVX1 port map( A => n3296, Y => n429);
   U402 : AOI22X1 port map( A0 => n430, A1 => n437, B0 => n3295, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248800_128249024_128249192, Y 
                           => n3296);
   U403 : OR3XL port map( A => output_signal_5_port, B => output_signal_6_port,
                           C => n3779, Y => n3777);
   U404 : XOR2X1 port map( A => n421, B => n3297, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128262496_128126088_128126312);
   U405 : XOR2X1 port map( A => n478, B => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128222208_128247288_128247512, Y 
                           => n3287);
   U406 : XOR2X1 port map( A => n449, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128248464_128248632, Y 
                           => n3293);
   U407 : XOR2X1 port map( A => n415, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128126480_128126592, Y 
                           => n3315);
   U408 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248016_128248128, B 
                           => n464, Y => n3305);
   U409 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248464_128248632, B 
                           => n460, Y => n3307);
   U410 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248856_128248968_128249136, B 
                           => n448, Y => n3309);
   U411 : XOR2X1 port map( A => n437, B => n430, Y => n3295);
   U412 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128249360_128249472_128249640, B 
                           => n438, Y => n3311);
   U413 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128222880_128247624_128247848, B 
                           => n3289, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124744_128124968_128125136);
   U414 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128247960_128248184_128248352, B 
                           => n3291, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125080_128125304_128125472);
   U415 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248296_128248520_128248688, B 
                           => n3293, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125416_128125640_128125808);
   U416 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248800_128249024_128249192, B 
                           => n3295, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125752_128125976_128126144);
   U417 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219288_128219512);
   U418 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219120_128219344);
   U419 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n481, Y => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219624_128219848);
   U420 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n472, Y => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer5_128219792_128220016);
   U421 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219456_128219680);
   U422 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219288_128219512);
   U423 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128247680_128247792, B 
                           => n3287, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124632_128124800_128124912);
   U424 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n472, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128219792_128220016);
   U425 : INVX1 port map( A => n3288, Y => n464);
   U426 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
                           A1 => n478, B0 => n3287, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128247680_128247792, Y 
                           => n3288);
   U427 : INVX1 port map( A => n3294, Y => n438);
   U428 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128248464_128248632, 
                           A1 => n449, B0 => n3293, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248296_128248520_128248688, Y 
                           => n3294);
   U429 : INVX1 port map( A => n3316, Y => n414);
   U430 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128126480_128126592, 
                           A1 => n415, B0 => n3315, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128263168_128126424_128126648, Y 
                           => n3316);
   U431 : INVX1 port map( A => n3306, Y => n452);
   U432 : AOI22X1 port map( A0 => n464, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248016_128248128, 
                           B0 => n3305, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124744_128124968_128125136, Y 
                           => n3306);
   U433 : INVX1 port map( A => n3308, Y => n440);
   U434 : AOI22X1 port map( A0 => n460, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248464_128248632, 
                           B0 => n3307, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125080_128125304_128125472, Y 
                           => n3308);
   U435 : INVX1 port map( A => n3310, Y => n431);
   U436 : AOI22X1 port map( A0 => n448, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
                           B0 => n3309, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125416_128125640_128125808, Y 
                           => n3310);
   U437 : INVX1 port map( A => n3312, Y => n422);
   U438 : AOI22X1 port map( A0 => n438, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
                           B0 => n3311, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128125752_128125976_128126144, Y 
                           => n3312);
   U439 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128126816_128126928, 
                           A1 => n418, B0 => n3317, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126760_128237640_128237808, Y 
                           => n3318);
   U440 : XOR2X1 port map( A => n3302, B => n29, Y => n3319);
   U441 : NAND2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => n29);
   U442 : AOI22X1 port map( A0 => n409, A1 => n412, B0 => n3301, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262664_128262888_128263056, Y 
                           => n3302);
   U443 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_5_port);
   U444 : XOR2X1 port map( A => n418, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128126816_128126928, Y 
                           => n3317);
   U445 : XOR2X1 port map( A => n412, B => n409, Y => n3301);
   U446 : OR3XL port map( A => output_previous_1_11_port, B => 
                           output_previous_1_12_port, C => n3788, Y => n3786);
   U447 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128126480_128126592);
   U448 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128126816_128126928);
   U449 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126816_128126928);
   U450 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128237920_128238088);
   U451 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126480_128126592);
   U452 : XOR2X1 port map( A => n425, B => n3299, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128263168_128126424_128126648);
   U453 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262664_128262888_128263056, B 
                           => n3301, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128126760_128237640_128237808);
   U454 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198080_128198192_128198360, B 
                           => n3279, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263224_128263392_128263504);
   U455 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224952_128225120_128225232, B 
                           => n3271, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128249696_128249808_128262328);
   U456 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197520_128197632_128197800, B 
                           => n3275, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262720_128262832_128263000);
   U457 : XNOR2X1 port map( A => n4000, B => n463, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_9_port);
   U458 : NOR3X1 port map( A => output_previous_1_13_port, B => 
                           output_previous_1_14_port, C => n3786, Y => n3785);
   U459 : NOR2BX1 port map( AN => n3785, B => output_previous_1_15_port, Y => 
                           n3784);
   U460 : INVX1 port map( A => output_previous_1_9_port, Y => n1210);
   U461 : XOR2X1 port map( A => n897, B => n2829, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128262496_128126088_128126312);
   U462 : XOR2X1 port map( A => n1056, B => n3063, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128262496_128126088_128126312);
   U463 : XOR2X1 port map( A => n579, B => n3531, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128262496_128126088_128126312);
   U464 : XOR2X1 port map( A => n738, B => n2595, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128262496_128126088_128126312);
   U465 : XOR2X1 port map( A => n913, B => n906, Y => n2827);
   U466 : XOR2X1 port map( A => n1072, B => n1065, Y => n3061);
   U467 : XOR2X1 port map( A => n595, B => n588, Y => n3529);
   U468 : XOR2X1 port map( A => n754, B => n747, Y => n2593);
   U469 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248800_128249024_128249192, B 
                           => n2827, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125752_128125976_128126144);
   U470 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248800_128249024_128249192, B 
                           => n2593, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125752_128125976_128126144);
   U471 : BUFX3 port map( A => n873, Y => n124);
   U472 : BUFX3 port map( A => n1032, Y => n128);
   U473 : BUFX3 port map( A => n555, Y => n116);
   U474 : BUFX3 port map( A => n714, Y => n120);
   U475 : INVX1 port map( A => n2828, Y => n905);
   U476 : AOI22X1 port map( A0 => n906, A1 => n913, B0 => n2827, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248800_128249024_128249192, Y 
                           => n2828);
   U477 : INVX1 port map( A => n3062, Y => n1064);
   U478 : AOI22X1 port map( A0 => n1065, A1 => n1072, B0 => n3061, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248800_128249024_128249192, Y 
                           => n3062);
   U479 : INVX1 port map( A => n3530, Y => n587);
   U480 : AOI22X1 port map( A0 => n588, A1 => n595, B0 => n3529, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248800_128249024_128249192, Y 
                           => n3530);
   U481 : INVX1 port map( A => n2594, Y => n746);
   U482 : AOI22X1 port map( A0 => n747, A1 => n754, B0 => n2593, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248800_128249024_128249192, Y 
                           => n2594);
   U483 : BUFX3 port map( A => n873, Y => n123);
   U484 : BUFX3 port map( A => n1032, Y => n127);
   U485 : BUFX3 port map( A => n555, Y => n115);
   U486 : BUFX3 port map( A => n714, Y => n119);
   U487 : NOR3X1 port map( A => n2311, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_8, C
                           => n3713, Y => n3711);
   U488 : NOR3X1 port map( A => n2332, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_8, C
                           => n3761, Y => n3759);
   U489 : NOR3X1 port map( A => n2374, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_8, 
                           C => n3857, Y => n3855);
   U490 : NOR3X1 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn47
                           , B => 
                           input_times_b0_mul_componentxunsigned_output_8, C =>
                           n3665, Y => n3663);
   U491 : INVX1 port map( A => n2826, Y => n914);
   U492 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128248464_128248632, 
                           A1 => n926, B0 => n2825, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248296_128248520_128248688, Y 
                           => n2826);
   U493 : INVX1 port map( A => n2592, Y => n755);
   U494 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128248464_128248632, 
                           A1 => n767, B0 => n2591, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248296_128248520_128248688, Y 
                           => n2592);
   U495 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128126816_128126928, 
                           A1 => n894, B0 => n2849, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126760_128237640_128237808, Y 
                           => n2850);
   U496 : INVX1 port map( A => n3082, Y => n1049);
   U497 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128126480_128126592, 
                           A1 => n1050, B0 => n3081, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128263168_128126424_128126648, Y 
                           => n3082);
   U498 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128126816_128126928, 
                           A1 => n1053, B0 => n3083, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126760_128237640_128237808, Y 
                           => n3084);
   U499 : INVX1 port map( A => n3550, Y => n572);
   U500 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128126480_128126592, 
                           A1 => n573, B0 => n3549, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128263168_128126424_128126648, Y 
                           => n3550);
   U501 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128126816_128126928, 
                           A1 => n576, B0 => n3551, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126760_128237640_128237808, Y 
                           => n3552);
   U502 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128126816_128126928, 
                           A1 => n735, B0 => n2615, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126760_128237640_128237808, Y 
                           => n2616);
   U503 : XOR2X1 port map( A => n955, B => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128222208_128247288_128247512, Y 
                           => n2819);
   U504 : XOR2X1 port map( A => n1114, B => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128222208_128247288_128247512, Y 
                           => n3053);
   U505 : XOR2X1 port map( A => n637, B => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128222208_128247288_128247512, Y 
                           => n3521);
   U506 : XOR2X1 port map( A => n796, B => 
                           input_times_b0_mul_componentxUMxsum_layer3_128222208_128247288_128247512, Y 
                           => n2585);
   U507 : XOR2X1 port map( A => n926, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128248464_128248632, Y 
                           => n2825);
   U508 : XOR2X1 port map( A => n1085, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128248464_128248632, Y 
                           => n3059);
   U509 : XOR2X1 port map( A => n608, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128248464_128248632, Y 
                           => n3527);
   U510 : XOR2X1 port map( A => n767, B => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128248464_128248632, Y 
                           => n2591);
   U511 : XOR2X1 port map( A => n891, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128126480_128126592, Y 
                           => n2847);
   U512 : XOR2X1 port map( A => n894, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128126816_128126928, Y 
                           => n2849);
   U513 : XOR2X1 port map( A => n1050, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128126480_128126592, Y 
                           => n3081);
   U514 : XOR2X1 port map( A => n1053, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128126816_128126928, Y 
                           => n3083);
   U515 : XOR2X1 port map( A => n573, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128126480_128126592, Y 
                           => n3549);
   U516 : XOR2X1 port map( A => n576, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128126816_128126928, Y 
                           => n3551);
   U517 : XOR2X1 port map( A => n732, B => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128126480_128126592, Y 
                           => n2613);
   U518 : XOR2X1 port map( A => n735, B => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128126816_128126928, Y 
                           => n2615);
   U519 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248016_128248128, B 
                           => n941, Y => n2837);
   U520 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248016_128248128, B 
                           => n1100, Y => n3071);
   U521 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248016_128248128, B 
                           => n623, Y => n3539);
   U522 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248016_128248128, B 
                           => n782, Y => n2603);
   U523 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248464_128248632, B 
                           => n937, Y => n2839);
   U524 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248464_128248632, B 
                           => n1096, Y => n3073);
   U525 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248464_128248632, B 
                           => n619, Y => n3541);
   U526 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248464_128248632, B 
                           => n778, Y => n2605);
   U527 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248856_128248968_128249136, B 
                           => n925, Y => n2841);
   U528 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248856_128248968_128249136, B 
                           => n1084, Y => n3075);
   U529 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248856_128248968_128249136, B 
                           => n607, Y => n3543);
   U530 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248856_128248968_128249136, B 
                           => n766, Y => n2607);
   U531 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128249360_128249472_128249640, B 
                           => n914, Y => n2843);
   U532 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128249360_128249472_128249640, B 
                           => n1073, Y => n3077);
   U533 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128249360_128249472_128249640, B 
                           => n596, Y => n3545);
   U534 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128249360_128249472_128249640, B 
                           => n755, Y => n2609);
   U535 : XOR2X1 port map( A => n888, B => n885, Y => n2833);
   U536 : XOR2X1 port map( A => n1047, B => n1044, Y => n3067);
   U537 : XOR2X1 port map( A => n570, B => n567, Y => n3535);
   U538 : XOR2X1 port map( A => n729, B => n726, Y => n2599);
   U539 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128126480_128126592);
   U540 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128126816_128126928);
   U541 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128126480_128126592);
   U542 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128126816_128126928);
   U543 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128126480_128126592);
   U544 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128126816_128126928);
   U545 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128126480_128126592);
   U546 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128126816_128126928);
   U547 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126816_128126928);
   U548 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126816_128126928);
   U549 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126816_128126928);
   U550 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262720_128262832_128263000, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262216_128262384_128262552, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126816_128126928);
   U551 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128222880_128247624_128247848, B 
                           => n2821, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124744_128124968_128125136);
   U552 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128222880_128247624_128247848, B 
                           => n3055, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124744_128124968_128125136);
   U553 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128222880_128247624_128247848, B 
                           => n3523, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124744_128124968_128125136);
   U554 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128222880_128247624_128247848, B 
                           => n2587, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124744_128124968_128125136);
   U555 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128247960_128248184_128248352, B 
                           => n2823, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125080_128125304_128125472);
   U556 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128247960_128248184_128248352, B 
                           => n3057, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125080_128125304_128125472);
   U557 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128247960_128248184_128248352, B 
                           => n3525, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125080_128125304_128125472);
   U558 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128247960_128248184_128248352, B 
                           => n2589, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125080_128125304_128125472);
   U559 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248296_128248520_128248688, B 
                           => n2825, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125416_128125640_128125808);
   U560 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248296_128248520_128248688, B 
                           => n3059, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125416_128125640_128125808);
   U561 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248296_128248520_128248688, B 
                           => n3527, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125416_128125640_128125808);
   U562 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248296_128248520_128248688, B 
                           => n2591, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125416_128125640_128125808);
   U563 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248800_128249024_128249192, B 
                           => n3061, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125752_128125976_128126144);
   U564 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248800_128249024_128249192, B 
                           => n3529, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125752_128125976_128126144);
   U565 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126480_128126592);
   U566 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126480_128126592);
   U567 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126480_128126592);
   U568 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128249696_128249808_128262328, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128197128_128249304_128249528, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126480_128126592);
   U569 : XOR2X1 port map( A => n901, B => n2831, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128263168_128126424_128126648);
   U570 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262664_128262888_128263056, B 
                           => n2833, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128126760_128237640_128237808);
   U571 : XOR2X1 port map( A => n1060, B => n3065, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128263168_128126424_128126648);
   U572 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262664_128262888_128263056, B 
                           => n3067, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128126760_128237640_128237808);
   U573 : XOR2X1 port map( A => n583, B => n3533, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128263168_128126424_128126648);
   U574 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262664_128262888_128263056, B 
                           => n3535, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128126760_128237640_128237808);
   U575 : XOR2X1 port map( A => n742, B => n2597, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128263168_128126424_128126648);
   U576 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262664_128262888_128263056, B 
                           => n2599, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128126760_128237640_128237808);
   U577 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219456_128219680);
   U578 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219288_128219512);
   U579 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219456_128219680);
   U580 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219288_128219512);
   U581 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219456_128219680);
   U582 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219288_128219512);
   U583 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219456_128219680);
   U584 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219288_128219512);
   U585 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n958, Y => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219624_128219848);
   U586 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n1117, Y => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219624_128219848);
   U587 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n640, Y => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219624_128219848);
   U588 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n799, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219624_128219848);
   U589 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n949, Y => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219792_128220016);
   U590 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n1108, Y => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219792_128220016);
   U591 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n631, Y => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219792_128220016);
   U592 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n790, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219792_128220016);
   U593 : XOR2X1 port map( A => n2834, B => n30, Y => n2851);
   U594 : NAND2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => n30);
   U595 : AOI22X1 port map( A0 => n885, A1 => n888, B0 => n2833, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262664_128262888_128263056, Y 
                           => n2834);
   U596 : XOR2X1 port map( A => n3068, B => n31, Y => n3085);
   U597 : NAND2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => n31);
   U598 : AOI22X1 port map( A0 => n1044, A1 => n1047, B0 => n3067, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262664_128262888_128263056, Y 
                           => n3068);
   U599 : XOR2X1 port map( A => n3536, B => n32, Y => n3553);
   U600 : NAND2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => n32);
   U601 : AOI22X1 port map( A0 => n567, A1 => n570, B0 => n3535, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262664_128262888_128263056, Y 
                           => n3536);
   U602 : XOR2X1 port map( A => n2600, B => n33, Y => n2617);
   U603 : NAND2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => n33);
   U604 : AOI22X1 port map( A0 => n726, A1 => n729, B0 => n2599, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262664_128262888_128263056, Y 
                           => n2600);
   U605 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219456_128219680);
   U606 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219288_128219512);
   U607 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219456_128219680);
   U608 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219456_128219680);
   U609 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128247120_128124240_128124520, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128124072_128124296, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219456_128219680);
   U610 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219288_128219512);
   U611 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246952_128247176_128247344, B 
                           => n2817, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128247456_128124464_128124688);
   U612 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246616_128246840_128247008, B 
                           => n2815, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128247120_128124240_128124520);
   U613 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246952_128247176_128247344, B 
                           => n3051, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128247456_128124464_128124688);
   U614 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246616_128246840_128247008, B 
                           => n3049, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128247120_128124240_128124520);
   U615 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246952_128247176_128247344, B 
                           => n3519, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128247456_128124464_128124688);
   U616 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246616_128246840_128247008, B 
                           => n3517, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128247120_128124240_128124520);
   U617 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246952_128247176_128247344, B 
                           => n2583, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128247456_128124464_128124688);
   U618 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246616_128246840_128247008, B 
                           => n2581, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128247120_128124240_128124520);
   U619 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128247680_128247792, B 
                           => n2819, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124632_128124800_128124912);
   U620 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128247680_128247792, B 
                           => n3053, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124632_128124800_128124912);
   U621 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128247680_128247792, B 
                           => n3521, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124632_128124800_128124912);
   U622 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128247680_128247792, B 
                           => n2585, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124632_128124800_128124912);
   U623 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n958, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219624_128219848);
   U624 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n1117, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219624_128219848);
   U625 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n640, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219624_128219848);
   U626 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128247456_128124464_128124688, B 
                           => n799, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219624_128219848);
   U627 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n949, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128219792_128220016);
   U628 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n1108, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219792_128220016);
   U629 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n631, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219792_128220016);
   U630 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124632_128124800_128124912, B 
                           => n790, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128219792_128220016);
   U631 : INVX1 port map( A => n2820, Y => n941);
   U632 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
                           A1 => n955, B0 => n2819, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128247680_128247792, Y 
                           => n2820);
   U633 : INVX1 port map( A => n3054, Y => n1100);
   U634 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
                           A1 => n1114, B0 => n3053, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128247680_128247792, Y 
                           => n3054);
   U635 : INVX1 port map( A => n3522, Y => n623);
   U636 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
                           A1 => n637, B0 => n3521, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128247680_128247792, Y 
                           => n3522);
   U637 : INVX1 port map( A => n2586, Y => n782);
   U638 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128222208_128247288_128247512, 
                           A1 => n796, B0 => n2585, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128247680_128247792, Y 
                           => n2586);
   U639 : INVX1 port map( A => n3060, Y => n1073);
   U640 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128248464_128248632, 
                           A1 => n1085, B0 => n3059, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248296_128248520_128248688, Y 
                           => n3060);
   U641 : INVX1 port map( A => n3528, Y => n596);
   U642 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128248464_128248632, 
                           A1 => n608, B0 => n3527, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248296_128248520_128248688, Y 
                           => n3528);
   U643 : INVX1 port map( A => n2848, Y => n890);
   U644 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128126480_128126592, 
                           A1 => n891, B0 => n2847, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128263168_128126424_128126648, Y 
                           => n2848);
   U645 : INVX1 port map( A => n2614, Y => n731);
   U646 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128126480_128126592, 
                           A1 => n732, B0 => n2613, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128263168_128126424_128126648, Y 
                           => n2614);
   U647 : INVX1 port map( A => n2838, Y => n929);
   U648 : AOI22X1 port map( A0 => n941, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248016_128248128, 
                           B0 => n2837, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124744_128124968_128125136, Y 
                           => n2838);
   U649 : INVX1 port map( A => n3072, Y => n1088);
   U650 : AOI22X1 port map( A0 => n1100, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248016_128248128, 
                           B0 => n3071, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124744_128124968_128125136, Y 
                           => n3072);
   U651 : INVX1 port map( A => n3540, Y => n611);
   U652 : AOI22X1 port map( A0 => n623, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248016_128248128, 
                           B0 => n3539, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124744_128124968_128125136, Y 
                           => n3540);
   U653 : INVX1 port map( A => n2604, Y => n770);
   U654 : AOI22X1 port map( A0 => n782, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248016_128248128, 
                           B0 => n2603, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124744_128124968_128125136, Y 
                           => n2604);
   U655 : INVX1 port map( A => n2840, Y => n916);
   U656 : AOI22X1 port map( A0 => n937, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248464_128248632, 
                           B0 => n2839, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125080_128125304_128125472, Y 
                           => n2840);
   U657 : INVX1 port map( A => n3074, Y => n1075);
   U658 : AOI22X1 port map( A0 => n1096, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248464_128248632, 
                           B0 => n3073, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125080_128125304_128125472, Y 
                           => n3074);
   U659 : INVX1 port map( A => n3542, Y => n598);
   U660 : AOI22X1 port map( A0 => n619, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248464_128248632, 
                           B0 => n3541, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125080_128125304_128125472, Y 
                           => n3542);
   U661 : INVX1 port map( A => n2606, Y => n757);
   U662 : AOI22X1 port map( A0 => n778, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248464_128248632, 
                           B0 => n2605, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125080_128125304_128125472, Y 
                           => n2606);
   U663 : INVX1 port map( A => n2842, Y => n907);
   U664 : AOI22X1 port map( A0 => n925, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
                           B0 => n2841, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125416_128125640_128125808, Y 
                           => n2842);
   U665 : INVX1 port map( A => n3076, Y => n1066);
   U666 : AOI22X1 port map( A0 => n1084, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
                           B0 => n3075, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125416_128125640_128125808, Y 
                           => n3076);
   U667 : INVX1 port map( A => n3544, Y => n589);
   U668 : AOI22X1 port map( A0 => n607, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
                           B0 => n3543, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125416_128125640_128125808, Y 
                           => n3544);
   U669 : INVX1 port map( A => n2608, Y => n748);
   U670 : AOI22X1 port map( A0 => n766, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248856_128248968_128249136, 
                           B0 => n2607, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125416_128125640_128125808, Y 
                           => n2608);
   U671 : INVX1 port map( A => n2844, Y => n898);
   U672 : AOI22X1 port map( A0 => n914, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
                           B0 => n2843, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128125752_128125976_128126144, Y 
                           => n2844);
   U673 : INVX1 port map( A => n3078, Y => n1057);
   U674 : AOI22X1 port map( A0 => n1073, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
                           B0 => n3077, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128125752_128125976_128126144, Y 
                           => n3078);
   U675 : INVX1 port map( A => n3546, Y => n580);
   U676 : AOI22X1 port map( A0 => n596, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
                           B0 => n3545, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128125752_128125976_128126144, Y 
                           => n3546);
   U677 : INVX1 port map( A => n2610, Y => n739);
   U678 : AOI22X1 port map( A0 => n755, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128249360_128249472_128249640, 
                           B0 => n2609, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer4_128125752_128125976_128126144, Y 
                           => n2610);
   U679 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_5_port);
   U680 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_5_port);
   U681 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_5_port);
   U682 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_5_port)
                           ;
   U683 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128237920_128238088);
   U684 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128237920_128238088);
   U685 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128237920_128238088);
   U686 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263672_128263840, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263224_128263392_128263504, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer4_128237920_128238088);
   U687 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer5_128219120_128219344);
   U688 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer5_128219120_128219344);
   U689 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer5_128219120_128219344);
   U690 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128123904_128124128, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128123792_128123960, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer5_128219120_128219344);
   U691 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128219288_128219512);
   U692 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124072_128124296, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128123904_128124128, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128219288_128219512);
   U693 : XNOR2X1 port map( A => n3914, B => n940, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_9_port);
   U694 : XNOR2X1 port map( A => n3957, B => n1099, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_9_port);
   U695 : XNOR2X1 port map( A => n4043, B => n622, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_9_port);
   U696 : XNOR2X1 port map( A => n3871, B => n781, Y => 
                           input_times_b0_div_componentxinput_A_inverted_9_port
                           );
   U697 : NAND3X1 port map( A => output_previous_1_11_port, B => 
                           output_previous_1_10_port, C => 
                           output_previous_1_12_port, Y => output_contracterxn5
                           );
   U698 : OR3XL port map( A => output_previous_1_12_port, B => 
                           output_previous_1_13_port, C => 
                           output_previous_1_14_port, Y => output_contracterxn8
                           );
   U699 : INVX1 port map( A => n3250, Y => n489);
   U700 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
                           A1 => n497, B0 => n3249, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827304_127827416, Y 
                           => n3250);
   U701 : XOR2X1 port map( A => n497, B => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127731808_127826912_127827136, Y 
                           => n3249);
   U702 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827752_127827920, B 
                           => n489, Y => n3283);
   U703 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221424_128221536_128221704, B 
                           => n482, Y => n3285);
   U704 : INVX1 port map( A => n232, Y => n398);
   U705 : BUFX3 port map( A => n1203, Y => n134);
   U706 : INVX1 port map( A => n3284, Y => n481);
   U707 : AOI22X1 port map( A0 => n489, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827752_127827920, 
                           B0 => n3283, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246616_128246840_128247008, Y 
                           => n3284);
   U708 : BUFX3 port map( A => n1203, Y => n133);
   U709 : NOR3X1 port map( A => n480, B => n473, C => n4001, Y => n4000);
   U710 : NOR3X1 port map( A => n423, B => n417, C => n4008, Y => n4007);
   U711 : INVX1 port map( A => n3254, Y => n478);
   U712 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127827752_127827920, 
                           A1 => n483, B0 => n3253, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827584_127827808_128221256, Y 
                           => n3254);
   U713 : INVX1 port map( A => n3260, Y => n449);
   U714 : AOI22X1 port map( A0 => n451, A1 => n457, B0 => n3259, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222376_128222600_128222768, Y 
                           => n3260);
   U715 : INVX1 port map( A => n3262, Y => n437);
   U716 : AOI22X1 port map( A0 => n439, A1 => n447, B0 => n3261, B1 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_128223384_128223552, Y 
                           => n3262);
   U717 : NAND3BX1 port map( AN => n453, B => n4547, C => n4000, Y => n4009);
   U718 : NOR2BX1 port map( AN => n4007, B => n408, Y => n4006);
   U719 : OR3XL port map( A => output_signal_3_port, B => output_signal_4_port,
                           C => n3781, Y => n3779);
   U720 : XOR2X1 port map( A => n471, B => n3255, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128222208_128247288_128247512);
   U721 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831456_127845712_127847616, B 
                           => n3215, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223440_128223608_128223776);
   U722 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673568_127675472_127730688, B 
                           => n3221, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224280_128224448_128224560);
   U723 : XOR2X1 port map( A => n483, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127827752_127827920, Y 
                           => n3253);
   U724 : XOR2X1 port map( A => n470, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128247680_128247792, Y 
                           => n3289);
   U725 : XOR2X1 port map( A => n459, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128248016_128248128, Y 
                           => n3291);
   U726 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127715424_128223048_128223272, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223440_128223608_128223776, Y 
                           => n3263);
   U727 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223720_128223944_128224168, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224280_128224448_128224560, Y 
                           => n3267);
   U728 : XOR2X1 port map( A => n457, B => n451, Y => n3259);
   U729 : XOR2X1 port map( A => n447, B => n439, Y => n3261);
   U730 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128196792_128196960_128197184, B 
                           => n433, Y => n3297);
   U731 : OR3XL port map( A => n441, B => n432, C => n4009, Y => n4008);
   U732 : OR3XL port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_5_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_6_port, C 
                           => n3811, Y => n3809);
   U733 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128247680_128247792);
   U734 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128248016_128248128);
   U735 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128248464_128248632);
   U736 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248016_128248128);
   U737 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223888_128224112_128224056, B 
                           => n3263, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248856_128248968_128249136);
   U738 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827248_127827472_127827640, B 
                           => n3251, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246616_128246840_128247008);
   U739 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827584_127827808_128221256, B 
                           => n3253, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246952_128247176_128247344);
   U740 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128247680_128247792);
   U741 : XOR2X1 port map( A => n461, B => n3257, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128222880_128247624_128247848);
   U742 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222376_128222600_128222768, B 
                           => n3259, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128247960_128248184_128248352);
   U743 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_128223384_128223552, B 
                           => n3261, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248296_128248520_128248688);
   U744 : XOR2X1 port map( A => n456, B => n3265, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248800_128249024_128249192);
   U745 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128246000_128246168);
   U746 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128123904_128124128);
   U747 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128123792_128123960);
   U748 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n496, Y => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer4_128124072_128124296);
   U749 : NAND2BX1 port map( AN => n401, B => n4006, Y => n4005);
   U750 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128123904_128124128);
   U751 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827304_127827416, B 
                           => n3249, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246504_128246672_128246784);
   U752 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127826576_127826800_127826968, B 
                           => n3247, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_127827080_128246280_128246560);
   U753 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n496, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128124072_128124296);
   U754 : INVX1 port map( A => n3290, Y => n460);
   U755 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128247680_128247792, 
                           A1 => n470, B0 => n3289, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128222880_128247624_128247848, Y 
                           => n3290);
   U756 : INVX1 port map( A => n3292, Y => n448);
   U757 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128248016_128248128, 
                           A1 => n459, B0 => n3291, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128247960_128248184_128248352, Y 
                           => n3292);
   U758 : INVX1 port map( A => n3264, Y => n430);
   U759 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
                           B0 => n3263, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223888_128224112_128224056, Y 
                           => n3264);
   U760 : XNOR2X1 port map( A => n4007, B => n408, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_15_port);
   U761 : XNOR2X1 port map( A => n4006, B => n401, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_16_port);
   U762 : XOR2X1 port map( A => n4008, B => n423, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_13_port);
   U763 : XNOR2X1 port map( A => n34, B => n417, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_14_port);
   U764 : NOR2X1 port map( A => n423, B => n4008, Y => n34);
   U765 : INVX1 port map( A => n3298, Y => n415);
   U766 : AOI22X1 port map( A0 => n433, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
                           B0 => n3297, B1 => n421, Y => n3298);
   U767 : INVX1 port map( A => n3268, Y => n421);
   U768 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
                           B0 => n3267, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224728_128224896_128225064, Y 
                           => n3268);
   U769 : INVX1 port map( A => n3286, Y => n472);
   U770 : AOI22X1 port map( A0 => n482, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
                           B0 => n3285, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246952_128247176_128247344, Y 
                           => n3286);
   U771 : INVX1 port map( A => n3300, Y => n418);
   U772 : AOI22X1 port map( A0 => n419, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198024_128197968, 
                           B0 => n3299, B1 => n425, Y => n3300);
   U773 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_3_port);
   U774 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_4_port);
   U775 : XOR2X1 port map( A => n454, B => n3237, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197464_128197688_128197856);
   U776 : XOR2X1 port map( A => n475, B => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224392_128224616_128224784, Y 
                           => n3271);
   U777 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831792_127846048_127847952, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673792_127675696_127730912, Y 
                           => n3235);
   U778 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127627392_128196680_128196848, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197016_128197240_128197352, Y 
                           => n3275);
   U779 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_128198024_128197968, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197464_128197688_128197856, Y 
                           => n3279);
   U780 : XOR2X1 port map( A => n428, B => n455, Y => n3219);
   U781 : XOR2X1 port map( A => n426, B => n446, Y => n3225);
   U782 : XOR2X1 port map( A => n444, B => n403, Y => n3237);
   U783 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198024_128197968, B 
                           => n419, Y => n3299);
   U784 : XOR2X1 port map( A => n424, B => n442, Y => n3273);
   U785 : OR3XL port map( A => n495, B => n488, C => n4002, Y => n4001);
   U786 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128248464_128248632);
   U787 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224728_128224896_128225064, B 
                           => n3267, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128249360_128249472_128249640);
   U788 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831680_127845936_127847840, B 
                           => n3227, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224952_128225120_128225232);
   U789 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732816_127722496_127724400, B 
                           => n3235, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197520_128197632_128197800);
   U790 : XOR2X1 port map( A => n406, B => n3277, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262664_128262888_128263056);
   U791 : OR3XL port map( A => n509, B => n503, C => n4003, Y => n4002);
   U792 : XOR2X1 port map( A => n420, B => n3269, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128197128_128249304_128249528);
   U793 : XOR2X1 port map( A => n413, B => n3273, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128262216_128262384_128262552);
   U794 : INVX1 port map( A => n4547, Y => n463);
   U795 : XOR2X1 port map( A => n3238, B => n3240, Y => n3281);
   U796 : AOI22X1 port map( A0 => n403, A1 => n444, B0 => n3237, B1 => n454, Y 
                           => n3238);
   U797 : INVX1 port map( A => n3276, Y => n409);
   U798 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
                           B0 => n3275, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197520_128197632_128197800, Y 
                           => n3276);
   U799 : XOR2X1 port map( A => n4009, B => n441, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_11_port);
   U800 : XNOR2X1 port map( A => n35, B => n432, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_12_port);
   U801 : NOR2X1 port map( A => n4009, B => n441, Y => n35);
   U802 : XOR2X1 port map( A => n4010, B => n453, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_10_port);
   U803 : NAND2X1 port map( A => n4000, B => n4547, Y => n4010);
   U804 : INVX1 port map( A => n3274, Y => n412);
   U805 : AOI22X1 port map( A0 => n442, A1 => n424, B0 => n3273, B1 => n413, Y 
                           => n3274);
   U806 : INVX1 port map( A => n3272, Y => n425);
   U807 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
                           A1 => n475, B0 => n3271, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224952_128225120_128225232, Y 
                           => n3272);
   U808 : XOR2X1 port map( A => n4177, B => n4178, Y => 
                           output_previous_1_13_port);
   U809 : XOR2X1 port map( A => n4181, B => n4182, Y => 
                           output_previous_1_11_port);
   U810 : XOR2X1 port map( A => n4176, B => n4175, Y => 
                           output_previous_1_14_port);
   U811 : XOR2X1 port map( A => n4154, B => n4155, Y => 
                           output_previous_1_8_port);
   U812 : XOR2X1 port map( A => n4184, B => n4183, Y => 
                           output_previous_1_10_port);
   U813 : XOR2X1 port map( A => n4180, B => n4179, Y => 
                           output_previous_1_12_port);
   U814 : XOR2X1 port map( A => n4152, B => n4153, Y => 
                           output_previous_1_9_port);
   U815 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_128198024_128197968, 
                           B0 => n3279, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198080_128198192_128198360, Y 
                           => n3280);
   U816 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673904_127675808_127731024, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732928_127722608_127724512, Y 
                           => n3241);
   U817 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831904_127846160_127848064, B 
                           => n3239, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198080_128198192_128198360);
   U818 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263672_128263840);
   U819 : XOR2X1 port map( A => n4001, B => n480, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_7_port);
   U820 : XNOR2X1 port map( A => n36, B => n473, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_8_port);
   U821 : NOR2X1 port map( A => n480, B => n4001, Y => n36);
   U822 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128263672_128263840, B 
                           => n3303, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128237752_128237976_128238144);
   U823 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128263672_128263840);
   U824 : XOR2X1 port map( A => n404, B => n402, Y => n3303);
   U825 : INVX1 port map( A => n3280, Y => n402);
   U826 : INVX1 port map( A => n3236, Y => n406);
   U827 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
                           B0 => n3235, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732816_127722496_127724400, Y 
                           => n3236);
   U828 : XOR2X1 port map( A => n4173, B => n4174, Y => 
                           output_previous_1_15_port);
   U829 : XOR2X1 port map( A => n4171, B => n1205, Y => 
                           output_previous_1_16_port);
   U830 : XOR2X1 port map( A => n4002, B => n495, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_5_port);
   U831 : XNOR2X1 port map( A => n37, B => n503, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_4_port);
   U832 : NOR2X1 port map( A => n509, B => n4003, Y => n37);
   U833 : XNOR2X1 port map( A => n38, B => n488, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_6_port);
   U834 : NOR2X1 port map( A => n495, B => n4002, Y => n38);
   U835 : BUFX3 port map( A => n80, Y => n114);
   U836 : BUFX3 port map( A => n80, Y => n113);
   U837 : XOR2X1 port map( A => n4003, B => n509, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_3_port);
   U838 : INVX1 port map( A => n2796, Y => n906);
   U839 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
                           B0 => n2795, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223888_128224112_128224056, Y 
                           => n2796);
   U840 : INVX1 port map( A => n2562, Y => n747);
   U841 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
                           B0 => n2561, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223888_128224112_128224056, Y 
                           => n2562);
   U842 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127715424_128223048_128223272, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223440_128223608_128223776, Y 
                           => n2795);
   U843 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127715424_128223048_128223272, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223440_128223608_128223776, Y 
                           => n3029);
   U844 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127715424_128223048_128223272, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223440_128223608_128223776, Y 
                           => n3497);
   U845 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127715424_128223048_128223272, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223440_128223608_128223776, Y 
                           => n2561);
   U846 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128196792_128196960_128197184, B 
                           => n909, Y => n2829);
   U847 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128196792_128196960_128197184, B 
                           => n1068, Y => n3063);
   U848 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128196792_128196960_128197184, B 
                           => n591, Y => n3531);
   U849 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128196792_128196960_128197184, B 
                           => n750, Y => n2595);
   U850 : INVX1 port map( A => n190, Y => n873);
   U851 : INVX1 port map( A => n211, Y => n1032);
   U852 : INVX1 port map( A => n253, Y => n555);
   U853 : INVX1 port map( A => n281, Y => n714);
   U854 : INVX1 port map( A => n3030, Y => n1065);
   U855 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
                           B0 => n3029, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223888_128224112_128224056, Y 
                           => n3030);
   U856 : INVX1 port map( A => n3498, Y => n588);
   U857 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223440_128223608_128223776, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127715424_128223048_128223272, 
                           B0 => n3497, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223888_128224112_128224056, Y 
                           => n3498);
   U858 : NOR3X1 port map( A => n899, B => n893, C => n3922, Y => n3921);
   U859 : NOR3X1 port map( A => n1058, B => n1052, C => n3965, Y => n3964);
   U860 : NOR3X1 port map( A => n581, B => n575, C => n4051, Y => n4050);
   U861 : NOR3X1 port map( A => n740, B => n734, C => n3879, Y => n3878);
   U862 : INVX1 port map( A => n2786, Y => n955);
   U863 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127827752_127827920, 
                           A1 => n960, B0 => n2785, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827584_127827808_128221256, Y 
                           => n2786);
   U864 : INVX1 port map( A => n3020, Y => n1114);
   U865 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127827752_127827920, 
                           A1 => n1119, B0 => n3019, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827584_127827808_128221256, Y 
                           => n3020);
   U866 : INVX1 port map( A => n3488, Y => n637);
   U867 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127827752_127827920, 
                           A1 => n642, B0 => n3487, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827584_127827808_128221256, Y 
                           => n3488);
   U868 : INVX1 port map( A => n2552, Y => n796);
   U869 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127827752_127827920, 
                           A1 => n801, B0 => n2551, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827584_127827808_128221256, Y 
                           => n2552);
   U870 : INVX1 port map( A => n2822, Y => n937);
   U871 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128247680_128247792, 
                           A1 => n947, B0 => n2821, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128222880_128247624_128247848, Y 
                           => n2822);
   U872 : INVX1 port map( A => n2588, Y => n778);
   U873 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128247680_128247792, 
                           A1 => n788, B0 => n2587, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128222880_128247624_128247848, Y 
                           => n2588);
   U874 : INVX1 port map( A => n2824, Y => n925);
   U875 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128248016_128248128, 
                           A1 => n936, B0 => n2823, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128247960_128248184_128248352, Y 
                           => n2824);
   U876 : INVX1 port map( A => n2794, Y => n913);
   U877 : AOI22X1 port map( A0 => n915, A1 => n924, B0 => n2793, B1 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_128223384_128223552, Y 
                           => n2794);
   U878 : INVX1 port map( A => n2590, Y => n766);
   U879 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128248016_128248128, 
                           A1 => n777, B0 => n2589, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128247960_128248184_128248352, Y 
                           => n2590);
   U880 : INVX1 port map( A => n2560, Y => n754);
   U881 : AOI22X1 port map( A0 => n756, A1 => n765, B0 => n2559, B1 => 
                           input_times_b0_mul_componentxUMxcarry_layer2_128223384_128223552, Y 
                           => n2560);
   U882 : INVX1 port map( A => n2808, Y => n885);
   U883 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
                           B0 => n2807, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197520_128197632_128197800, Y 
                           => n2808);
   U884 : INVX1 port map( A => n2574, Y => n726);
   U885 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
                           B0 => n2573, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197520_128197632_128197800, Y 
                           => n2574);
   U886 : INVX1 port map( A => n2830, Y => n891);
   U887 : AOI22X1 port map( A0 => n909, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
                           B0 => n2829, B1 => n897, Y => n2830);
   U888 : INVX1 port map( A => n2832, Y => n894);
   U889 : AOI22X1 port map( A0 => n895, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198024_128197968, 
                           B0 => n2831, B1 => n901, Y => n2832);
   U890 : INVX1 port map( A => n3040, Y => n1047);
   U891 : AOI22X1 port map( A0 => n1077, A1 => n1059, B0 => n3039, B1 => n1048,
                           Y => n3040);
   U892 : INVX1 port map( A => n3508, Y => n570);
   U893 : AOI22X1 port map( A0 => n600, A1 => n582, B0 => n3507, B1 => n571, Y 
                           => n3508);
   U894 : INVX1 port map( A => n2596, Y => n732);
   U895 : AOI22X1 port map( A0 => n750, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
                           B0 => n2595, B1 => n738, Y => n2596);
   U896 : INVX1 port map( A => n2598, Y => n735);
   U897 : AOI22X1 port map( A0 => n736, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198024_128197968, 
                           B0 => n2597, B1 => n742, Y => n2598);
   U898 : NAND3BX1 port map( AN => n930, B => n4441, C => n3914, Y => n3923);
   U899 : NAND3BX1 port map( AN => n1089, B => n4494, C => n3957, Y => n3966);
   U900 : NAND3BX1 port map( AN => n612, B => n4600, C => n4043, Y => n4052);
   U901 : NAND3BX1 port map( AN => n771, B => input_times_b0_mul_componentxn90,
                           C => n3871, Y => n3880);
   U902 : NOR2BX1 port map( AN => n3921, B => n884, Y => n3920);
   U903 : NOR2BX1 port map( AN => n3964, B => n1043, Y => n3963);
   U904 : NOR2BX1 port map( AN => n4050, B => n566, Y => n4049);
   U905 : NOR2BX1 port map( AN => n3878, B => n725, Y => n3877);
   U906 : XOR2X1 port map( A => n948, B => n2787, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128222208_128247288_128247512);
   U907 : XOR2X1 port map( A => n1107, B => n3021, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128222208_128247288_128247512);
   U908 : XOR2X1 port map( A => n630, B => n3489, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128222208_128247288_128247512);
   U909 : XOR2X1 port map( A => n789, B => n2553, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128222208_128247288_128247512);
   U910 : XOR2X1 port map( A => n974, B => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127731808_127826912_127827136, Y 
                           => n2781);
   U911 : XOR2X1 port map( A => n1133, B => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127731808_127826912_127827136, Y 
                           => n3015);
   U912 : XOR2X1 port map( A => n656, B => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127731808_127826912_127827136, Y 
                           => n3483);
   U913 : XOR2X1 port map( A => n815, B => 
                           input_times_b0_mul_componentxUMxsum_layer2_127731808_127826912_127827136, Y 
                           => n2547);
   U914 : XOR2X1 port map( A => n960, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127827752_127827920, Y 
                           => n2785);
   U915 : XOR2X1 port map( A => n1119, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127827752_127827920, Y 
                           => n3019);
   U916 : XOR2X1 port map( A => n642, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127827752_127827920, Y 
                           => n3487);
   U917 : XOR2X1 port map( A => n801, B => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127827752_127827920, Y 
                           => n2551);
   U918 : XOR2X1 port map( A => n947, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128247680_128247792, Y 
                           => n2821);
   U919 : XOR2X1 port map( A => n936, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128248016_128248128, Y 
                           => n2823);
   U920 : XOR2X1 port map( A => n1106, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128247680_128247792, Y 
                           => n3055);
   U921 : XOR2X1 port map( A => n1095, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128248016_128248128, Y 
                           => n3057);
   U922 : XOR2X1 port map( A => n629, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128247680_128247792, Y 
                           => n3523);
   U923 : XOR2X1 port map( A => n618, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128248016_128248128, Y 
                           => n3525);
   U924 : XOR2X1 port map( A => n788, B => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128247680_128247792, Y 
                           => n2587);
   U925 : XOR2X1 port map( A => n777, B => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128248016_128248128, Y 
                           => n2589);
   U926 : XOR2X1 port map( A => n952, B => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224392_128224616_128224784, Y 
                           => n2803);
   U927 : XOR2X1 port map( A => n1111, B => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224392_128224616_128224784, Y 
                           => n3037);
   U928 : XOR2X1 port map( A => n634, B => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224392_128224616_128224784, Y 
                           => n3505);
   U929 : XOR2X1 port map( A => n793, B => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224392_128224616_128224784, Y 
                           => n2569);
   U930 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223720_128223944_128224168, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224280_128224448_128224560, Y 
                           => n2799);
   U931 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223720_128223944_128224168, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224280_128224448_128224560, Y 
                           => n3033);
   U932 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223720_128223944_128224168, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224280_128224448_128224560, Y 
                           => n3501);
   U933 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223720_128223944_128224168, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224280_128224448_128224560, Y 
                           => n2565);
   U934 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127627392_128196680_128196848, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197016_128197240_128197352, Y 
                           => n2807);
   U935 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127627392_128196680_128196848, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197016_128197240_128197352, Y 
                           => n3041);
   U936 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127627392_128196680_128196848, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197016_128197240_128197352, Y 
                           => n3509);
   U937 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127627392_128196680_128196848, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197016_128197240_128197352, Y 
                           => n2573);
   U938 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827752_127827920, B 
                           => n966, Y => n2815);
   U939 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827752_127827920, B 
                           => n1125, Y => n3049);
   U940 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827752_127827920, B 
                           => n648, Y => n3517);
   U941 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827752_127827920, B 
                           => n807, Y => n2581);
   U942 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221424_128221536_128221704, B 
                           => n959, Y => n2817);
   U943 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221424_128221536_128221704, B 
                           => n1118, Y => n3051);
   U944 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221424_128221536_128221704, B 
                           => n641, Y => n3519);
   U945 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221424_128221536_128221704, B 
                           => n800, Y => n2583);
   U946 : XOR2X1 port map( A => n934, B => n928, Y => n2791);
   U947 : XOR2X1 port map( A => n1093, B => n1087, Y => n3025);
   U948 : XOR2X1 port map( A => n616, B => n610, Y => n3493);
   U949 : XOR2X1 port map( A => n775, B => n769, Y => n2557);
   U950 : XOR2X1 port map( A => n924, B => n915, Y => n2793);
   U951 : XOR2X1 port map( A => n1083, B => n1074, Y => n3027);
   U952 : XOR2X1 port map( A => n606, B => n597, Y => n3495);
   U953 : XOR2X1 port map( A => n765, B => n756, Y => n2559);
   U954 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198024_128197968, B 
                           => n895, Y => n2831);
   U955 : XOR2X1 port map( A => n900, B => n918, Y => n2805);
   U956 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198024_128197968, B 
                           => n1054, Y => n3065);
   U957 : XOR2X1 port map( A => n1059, B => n1077, Y => n3039);
   U958 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198024_128197968, B 
                           => n577, Y => n3533);
   U959 : XOR2X1 port map( A => n582, B => n600, Y => n3507);
   U960 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198024_128197968, B 
                           => n736, Y => n2597);
   U961 : XOR2X1 port map( A => n741, B => n759, Y => n2571);
   U962 : OR3XL port map( A => n917, B => n908, C => n3923, Y => n3922);
   U963 : OR3XL port map( A => n1076, B => n1067, C => n3966, Y => n3965);
   U964 : OR3XL port map( A => n599, B => n590, C => n4052, Y => n4051);
   U965 : OR3XL port map( A => n758, B => n749, C => n3880, Y => n3879);
   U966 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128248016_128248128);
   U967 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128247680_128247792);
   U968 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128248016_128248128);
   U969 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128247680_128247792);
   U970 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128248016_128248128);
   U971 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128247680_128247792);
   U972 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128248016_128248128);
   U973 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128247680_128247792);
   U974 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128248464_128248632);
   U975 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128248464_128248632);
   U976 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128248464_128248632);
   U977 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128248464_128248632);
   U978 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248464_128248632);
   U979 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248464_128248632);
   U980 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248464_128248632);
   U981 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223384_128223552, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222936_128223104_128223216, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248464_128248632);
   U982 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223888_128224112_128224056, B 
                           => n2795, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248856_128248968_128249136);
   U983 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223888_128224112_128224056, B 
                           => n3029, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248856_128248968_128249136);
   U984 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223888_128224112_128224056, B 
                           => n3497, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248856_128248968_128249136);
   U985 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223888_128224112_128224056, B 
                           => n2561, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248856_128248968_128249136);
   U986 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224728_128224896_128225064, B 
                           => n2799, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128249360_128249472_128249640);
   U987 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224728_128224896_128225064, B 
                           => n3033, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128249360_128249472_128249640);
   U988 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224728_128224896_128225064, B 
                           => n3501, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128249360_128249472_128249640);
   U989 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224728_128224896_128225064, B 
                           => n2565, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128249360_128249472_128249640);
   U990 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827248_127827472_127827640, B 
                           => n2783, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246616_128246840_128247008);
   U991 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827248_127827472_127827640, B 
                           => n3017, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246616_128246840_128247008);
   U992 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827248_127827472_127827640, B 
                           => n3485, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246616_128246840_128247008);
   U993 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827248_127827472_127827640, B 
                           => n2549, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246616_128246840_128247008);
   U994 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827584_127827808_128221256, B 
                           => n2785, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246952_128247176_128247344);
   U995 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827584_127827808_128221256, B 
                           => n3019, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246952_128247176_128247344);
   U996 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827584_127827808_128221256, B 
                           => n3487, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246952_128247176_128247344);
   U997 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827584_127827808_128221256, B 
                           => n2551, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246952_128247176_128247344);
   U998 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128247680_128247792);
   U999 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128247680_128247792);
   U1000 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128247680_128247792);
   U1001 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221760_128221928_128222040, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_127635584_128221368_128221592, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128247680_128247792);
   U1002 : XOR2X1 port map( A => n938, B => n2789, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128222880_128247624_128247848);
   U1003 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222376_128222600_128222768, B 
                           => n2791, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128247960_128248184_128248352);
   U1004 : XOR2X1 port map( A => n1097, B => n3023, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128222880_128247624_128247848);
   U1005 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222376_128222600_128222768, B 
                           => n3025, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128247960_128248184_128248352);
   U1006 : XOR2X1 port map( A => n620, B => n3491, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128222880_128247624_128247848);
   U1007 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222376_128222600_128222768, B 
                           => n3493, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128247960_128248184_128248352);
   U1008 : XOR2X1 port map( A => n779, B => n2555, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128222880_128247624_128247848);
   U1009 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222376_128222600_128222768, B 
                           => n2557, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128247960_128248184_128248352);
   U1010 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_128223384_128223552, B 
                           => n2793, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248296_128248520_128248688);
   U1011 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_128223384_128223552, B 
                           => n3027, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248296_128248520_128248688);
   U1012 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_128223384_128223552, B 
                           => n3495, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248296_128248520_128248688);
   U1013 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxcarry_layer2_128223384_128223552, B 
                           => n2559, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248296_128248520_128248688);
   U1014 : XOR2X1 port map( A => n933, B => n2797, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248800_128249024_128249192);
   U1015 : XOR2X1 port map( A => n1092, B => n3031, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248800_128249024_128249192);
   U1016 : XOR2X1 port map( A => n615, B => n3499, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248800_128249024_128249192);
   U1017 : XOR2X1 port map( A => n774, B => n2563, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248800_128249024_128249192);
   U1018 : XOR2X1 port map( A => n896, B => n2801, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128197128_128249304_128249528);
   U1019 : XOR2X1 port map( A => n889, B => n2805, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262216_128262384_128262552);
   U1020 : XOR2X1 port map( A => n1055, B => n3035, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128197128_128249304_128249528);
   U1021 : XOR2X1 port map( A => n1048, B => n3039, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262216_128262384_128262552);
   U1022 : XOR2X1 port map( A => n578, B => n3503, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128197128_128249304_128249528);
   U1023 : XOR2X1 port map( A => n571, B => n3507, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262216_128262384_128262552);
   U1024 : XOR2X1 port map( A => n737, B => n2567, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128197128_128249304_128249528);
   U1025 : XOR2X1 port map( A => n730, B => n2571, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262216_128262384_128262552);
   U1026 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128123904_128124128);
   U1027 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128123904_128124128);
   U1028 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128123904_128124128);
   U1029 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128123904_128124128);
   U1030 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n973, Y => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128124072_128124296);
   U1031 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n1132, Y => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128124072_128124296);
   U1032 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n655, Y => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128124072_128124296);
   U1033 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n814, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128124072_128124296);
   U1034 : NAND2BX1 port map( AN => n876, B => n3920, Y => n3919);
   U1035 : NAND2BX1 port map( AN => n1035, B => n3963, Y => n3962);
   U1036 : NAND2BX1 port map( AN => n558, B => n4049, Y => n4048);
   U1037 : NAND2BX1 port map( AN => n717, B => n3877, Y => n3876);
   U1038 : XOR2X1 port map( A => n875, B => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_17_port, Y 
                           => n2313);
   U1039 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128315744_128315968_128316136, B 
                           => n2856, Y => 
                           input_p1_times_b1_mul_componentxUMxsecond_vector_17_port);
   U1040 : INVX1 port map( A => n2855, Y => n875);
   U1041 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128237752_128237976_128238144, B 
                           => n2851, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer5_128315744_128315968_128316136);
   U1042 : XOR2X1 port map( A => n1034, B => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_17_port, Y 
                           => n2334);
   U1043 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128315744_128315968_128316136, B 
                           => n3090, Y => 
                           input_p2_times_b2_mul_componentxUMxsecond_vector_17_port);
   U1044 : INVX1 port map( A => n3089, Y => n1034);
   U1045 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128237752_128237976_128238144, B 
                           => n3085, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer5_128315744_128315968_128316136);
   U1046 : XOR2X1 port map( A => n557, B => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_17_port, Y 
                           => n2376);
   U1047 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128315744_128315968_128316136, B 
                           => n3558, Y => 
                           output_p2_times_a2_mul_componentxUMxsecond_vector_17_port);
   U1048 : INVX1 port map( A => n3557, Y => n557);
   U1049 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128237752_128237976_128238144, B 
                           => n3553, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer5_128315744_128315968_128316136);
   U1050 : XOR2X1 port map( A => n716, B => 
                           input_times_b0_mul_componentxUMxsecond_vector_17_port, Y 
                           => input_times_b0_mul_componentxUMxAdder_finalxn475)
                           ;
   U1051 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer5_128315744_128315968_128316136, B 
                           => n2622, Y => 
                           input_times_b0_mul_componentxUMxsecond_vector_17_port);
   U1052 : INVX1 port map( A => n2621, Y => n716);
   U1053 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128237752_128237976_128238144, B 
                           => n2617, Y => 
                           input_times_b0_mul_componentxUMxsum_layer5_128315744_128315968_128316136);
   U1054 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827304_127827416, B 
                           => n2781, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246504_128246672_128246784);
   U1055 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127826576_127826800_127826968, B 
                           => n2779, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_127827080_128246280_128246560);
   U1056 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827304_127827416, B 
                           => n3015, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246504_128246672_128246784);
   U1057 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127826576_127826800_127826968, B 
                           => n3013, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_127827080_128246280_128246560);
   U1058 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827304_127827416, B 
                           => n3483, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246504_128246672_128246784);
   U1059 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127826576_127826800_127826968, B 
                           => n3481, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_127827080_128246280_128246560);
   U1060 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827304_127827416, B 
                           => n2547, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246504_128246672_128246784);
   U1061 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127826576_127826800_127826968, B 
                           => n2545, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_127827080_128246280_128246560);
   U1062 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224952_128225120_128225232, B 
                           => n2803, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128249696_128249808_128262328);
   U1063 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197520_128197632_128197800, B 
                           => n2807, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262720_128262832_128263000);
   U1064 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224952_128225120_128225232, B 
                           => n3037, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128249696_128249808_128262328);
   U1065 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197520_128197632_128197800, B 
                           => n3041, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262720_128262832_128263000);
   U1066 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224952_128225120_128225232, B 
                           => n3505, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128249696_128249808_128262328);
   U1067 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197520_128197632_128197800, B 
                           => n3509, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262720_128262832_128263000);
   U1068 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224952_128225120_128225232, B 
                           => n2569, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128249696_128249808_128262328);
   U1069 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197520_128197632_128197800, B 
                           => n2573, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262720_128262832_128263000);
   U1070 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n973, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128124072_128124296);
   U1071 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n1132, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128124072_128124296);
   U1072 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n655, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128124072_128124296);
   U1073 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246504_128246672_128246784, B 
                           => n814, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128124072_128124296);
   U1074 : INVX1 port map( A => n2782, Y => n966);
   U1075 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
                           A1 => n974, B0 => n2781, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827304_127827416, Y 
                           => n2782);
   U1076 : INVX1 port map( A => n3016, Y => n1125);
   U1077 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
                           A1 => n1133, B0 => n3015, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827304_127827416, Y 
                           => n3016);
   U1078 : INVX1 port map( A => n3484, Y => n648);
   U1079 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
                           A1 => n656, B0 => n3483, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827304_127827416, Y 
                           => n3484);
   U1080 : INVX1 port map( A => n2548, Y => n807);
   U1081 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer2_127731808_127826912_127827136, 
                           A1 => n815, B0 => n2547, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827304_127827416, Y 
                           => n2548);
   U1082 : INVX1 port map( A => n3056, Y => n1096);
   U1083 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128247680_128247792, 
                           A1 => n1106, B0 => n3055, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128222880_128247624_128247848, Y 
                           => n3056);
   U1084 : INVX1 port map( A => n3524, Y => n619);
   U1085 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128247680_128247792, 
                           A1 => n629, B0 => n3523, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128222880_128247624_128247848, Y 
                           => n3524);
   U1086 : INVX1 port map( A => n3058, Y => n1084);
   U1087 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128248016_128248128, 
                           A1 => n1095, B0 => n3057, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128247960_128248184_128248352, Y 
                           => n3058);
   U1088 : INVX1 port map( A => n3526, Y => n607);
   U1089 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128248016_128248128, 
                           A1 => n618, B0 => n3525, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128247960_128248184_128248352, Y 
                           => n3526);
   U1090 : INVX1 port map( A => n3042, Y => n1044);
   U1091 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
                           B0 => n3041, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197520_128197632_128197800, Y 
                           => n3042);
   U1092 : INVX1 port map( A => n3510, Y => n567);
   U1093 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197016_128197240_128197352, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127627392_128196680_128196848, 
                           B0 => n3509, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197520_128197632_128197800, Y 
                           => n3510);
   U1094 : XNOR2X1 port map( A => n3921, B => n884, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_15_port);
   U1095 : XNOR2X1 port map( A => n3964, B => n1043, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_15_port);
   U1096 : XNOR2X1 port map( A => n4050, B => n566, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_15_port);
   U1097 : XNOR2X1 port map( A => n3878, B => n725, Y => 
                           input_times_b0_div_componentxinput_A_inverted_15_port);
   U1098 : XNOR2X1 port map( A => n3920, B => n876, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_16_port);
   U1099 : XNOR2X1 port map( A => n3963, B => n1035, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_16_port);
   U1100 : XNOR2X1 port map( A => n4049, B => n558, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_16_port);
   U1101 : XNOR2X1 port map( A => n3877, B => n717, Y => 
                           input_times_b0_div_componentxinput_A_inverted_16_port);
   U1102 : XNOR2X1 port map( A => n39, B => n893, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_14_port);
   U1103 : NOR2X1 port map( A => n899, B => n3922, Y => n39);
   U1104 : XNOR2X1 port map( A => n40, B => n1052, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_14_port);
   U1105 : NOR2X1 port map( A => n1058, B => n3965, Y => n40);
   U1106 : XNOR2X1 port map( A => n41, B => n575, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_14_port);
   U1107 : NOR2X1 port map( A => n581, B => n4051, Y => n41);
   U1108 : XNOR2X1 port map( A => n42, B => n734, Y => 
                           input_times_b0_div_componentxinput_A_inverted_14_port);
   U1109 : NOR2X1 port map( A => n740, B => n3879, Y => n42);
   U1110 : INVX1 port map( A => n2792, Y => n926);
   U1111 : AOI22X1 port map( A0 => n928, A1 => n934, B0 => n2791, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222376_128222600_128222768, Y 
                           => n2792);
   U1112 : INVX1 port map( A => n3026, Y => n1085);
   U1113 : AOI22X1 port map( A0 => n1087, A1 => n1093, B0 => n3025, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222376_128222600_128222768, Y 
                           => n3026);
   U1114 : INVX1 port map( A => n3494, Y => n608);
   U1115 : AOI22X1 port map( A0 => n610, A1 => n616, B0 => n3493, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222376_128222600_128222768, Y 
                           => n3494);
   U1116 : INVX1 port map( A => n2558, Y => n767);
   U1117 : AOI22X1 port map( A0 => n769, A1 => n775, B0 => n2557, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222376_128222600_128222768, Y 
                           => n2558);
   U1118 : INVX1 port map( A => n3028, Y => n1072);
   U1119 : AOI22X1 port map( A0 => n1074, A1 => n1083, B0 => n3027, B1 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_128223384_128223552, Y 
                           => n3028);
   U1120 : INVX1 port map( A => n3496, Y => n595);
   U1121 : AOI22X1 port map( A0 => n597, A1 => n606, B0 => n3495, B1 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_128223384_128223552, Y 
                           => n3496);
   U1122 : INVX1 port map( A => n2806, Y => n888);
   U1123 : AOI22X1 port map( A0 => n918, A1 => n900, B0 => n2805, B1 => n889, Y
                           => n2806);
   U1124 : INVX1 port map( A => n3064, Y => n1050);
   U1125 : AOI22X1 port map( A0 => n1068, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
                           B0 => n3063, B1 => n1056, Y => n3064);
   U1126 : INVX1 port map( A => n3066, Y => n1053);
   U1127 : AOI22X1 port map( A0 => n1054, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198024_128197968, 
                           B0 => n3065, B1 => n1060, Y => n3066);
   U1128 : INVX1 port map( A => n3532, Y => n573);
   U1129 : AOI22X1 port map( A0 => n591, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128196792_128196960_128197184, 
                           B0 => n3531, B1 => n579, Y => n3532);
   U1130 : INVX1 port map( A => n3534, Y => n576);
   U1131 : AOI22X1 port map( A0 => n577, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198024_128197968, 
                           B0 => n3533, B1 => n583, Y => n3534);
   U1132 : INVX1 port map( A => n2572, Y => n729);
   U1133 : AOI22X1 port map( A0 => n759, A1 => n741, B0 => n2571, B1 => n730, Y
                           => n2572);
   U1134 : INVX1 port map( A => n2800, Y => n897);
   U1135 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
                           B0 => n2799, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224728_128224896_128225064, Y 
                           => n2800);
   U1136 : INVX1 port map( A => n2804, Y => n901);
   U1137 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
                           A1 => n952, B0 => n2803, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224952_128225120_128225232, Y 
                           => n2804);
   U1138 : INVX1 port map( A => n3034, Y => n1056);
   U1139 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
                           B0 => n3033, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224728_128224896_128225064, Y 
                           => n3034);
   U1140 : INVX1 port map( A => n3038, Y => n1060);
   U1141 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
                           A1 => n1111, B0 => n3037, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224952_128225120_128225232, Y 
                           => n3038);
   U1142 : INVX1 port map( A => n3502, Y => n579);
   U1143 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
                           B0 => n3501, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224728_128224896_128225064, Y 
                           => n3502);
   U1144 : INVX1 port map( A => n3506, Y => n583);
   U1145 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
                           A1 => n634, B0 => n3505, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224952_128225120_128225232, Y 
                           => n3506);
   U1146 : INVX1 port map( A => n2566, Y => n738);
   U1147 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224280_128224448_128224560, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223720_128223944_128224168, 
                           B0 => n2565, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224728_128224896_128225064, Y 
                           => n2566);
   U1148 : INVX1 port map( A => n2570, Y => n742);
   U1149 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224392_128224616_128224784, 
                           A1 => n793, B0 => n2569, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224952_128225120_128225232, Y 
                           => n2570);
   U1150 : INVX1 port map( A => n2816, Y => n958);
   U1151 : AOI22X1 port map( A0 => n966, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827752_127827920, 
                           B0 => n2815, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246616_128246840_128247008, Y 
                           => n2816);
   U1152 : INVX1 port map( A => n3050, Y => n1117);
   U1153 : AOI22X1 port map( A0 => n1125, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827752_127827920, 
                           B0 => n3049, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246616_128246840_128247008, Y 
                           => n3050);
   U1154 : INVX1 port map( A => n3518, Y => n640);
   U1155 : AOI22X1 port map( A0 => n648, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827752_127827920, 
                           B0 => n3517, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246616_128246840_128247008, Y 
                           => n3518);
   U1156 : INVX1 port map( A => n2582, Y => n799);
   U1157 : AOI22X1 port map( A0 => n807, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827752_127827920, 
                           B0 => n2581, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246616_128246840_128247008, Y 
                           => n2582);
   U1158 : INVX1 port map( A => n2818, Y => n949);
   U1159 : AOI22X1 port map( A0 => n959, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
                           B0 => n2817, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246952_128247176_128247344, Y 
                           => n2818);
   U1160 : INVX1 port map( A => n3052, Y => n1108);
   U1161 : AOI22X1 port map( A0 => n1118, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
                           B0 => n3051, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246952_128247176_128247344, Y 
                           => n3052);
   U1162 : INVX1 port map( A => n3520, Y => n631);
   U1163 : AOI22X1 port map( A0 => n641, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
                           B0 => n3519, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246952_128247176_128247344, Y 
                           => n3520);
   U1164 : INVX1 port map( A => n2584, Y => n790);
   U1165 : AOI22X1 port map( A0 => n800, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221424_128221536_128221704, 
                           B0 => n2583, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246952_128247176_128247344, Y 
                           => n2584);
   U1166 : NOR3X1 port map( A => n957, B => n950, C => n3915, Y => n3914);
   U1167 : NOR3X1 port map( A => n1116, B => n1109, C => n3958, Y => n3957);
   U1168 : NOR3X1 port map( A => n639, B => n632, C => n4044, Y => n4043);
   U1169 : NOR3X1 port map( A => n798, B => n791, C => n3872, Y => n3871);
   U1170 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_4_port);
   U1171 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_4_port);
   U1172 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_4_port);
   U1173 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_4_port)
                           ;
   U1174 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_128198024_128197968, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197464_128197688_128197856, Y 
                           => n2811);
   U1175 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_128198024_128197968, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197464_128197688_128197856, Y 
                           => n3045);
   U1176 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_128198024_128197968, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197464_128197688_128197856, Y 
                           => n3513);
   U1177 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxcarry_layer2_128198024_128197968, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197464_128197688_128197856, Y 
                           => n2577);
   U1178 : OR3XL port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_5_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_6_port, C 
                           => n3715, Y => n3713);
   U1179 : OR3XL port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_5_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_6_port, C 
                           => n3763, Y => n3761);
   U1180 : OR3XL port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_5_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_6_port, C 
                           => n3859, Y => n3857);
   U1181 : OR3XL port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_5_port,
                           B => 
                           input_times_b0_mul_componentxUMxfirst_vector_6_port,
                           C => n3667, Y => n3665);
   U1182 : OR3XL port map( A => n972, B => n965, C => n3916, Y => n3915);
   U1183 : OR3XL port map( A => n1131, B => n1124, C => n3959, Y => n3958);
   U1184 : OR3XL port map( A => n654, B => n647, C => n4045, Y => n4044);
   U1185 : OR3XL port map( A => n813, B => n806, C => n3873, Y => n3872);
   U1186 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128248016_128248128);
   U1187 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128248016_128248128);
   U1188 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128248016_128248128);
   U1189 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222432_128222544_128222712, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221872_128222096_128222264, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128248016_128248128);
   U1190 : XOR2X1 port map( A => n882, B => n2809, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128262664_128262888_128263056);
   U1191 : XOR2X1 port map( A => n1041, B => n3043, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128262664_128262888_128263056);
   U1192 : XOR2X1 port map( A => n564, B => n3511, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128262664_128262888_128263056);
   U1193 : XOR2X1 port map( A => n723, B => n2575, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128262664_128262888_128263056);
   U1194 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198080_128198192_128198360, B 
                           => n2811, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263224_128263392_128263504);
   U1195 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198080_128198192_128198360, B 
                           => n3045, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263224_128263392_128263504);
   U1196 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198080_128198192_128198360, B 
                           => n3513, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263224_128263392_128263504);
   U1197 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198080_128198192_128198360, B 
                           => n2577, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263224_128263392_128263504);
   U1198 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128246000_128246168);
   U1199 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128246000_128246168);
   U1200 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128246000_128246168);
   U1201 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128246000_128246168);
   U1202 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer4_128123792_128123960);
   U1203 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer4_128123792_128123960);
   U1204 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer4_128123792_128123960);
   U1205 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246112_128246336, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128246000_128246168, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer4_128123792_128123960);
   U1206 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128123904_128124128);
   U1207 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128123904_128124128);
   U1208 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128123904_128124128);
   U1209 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_127827080_128246280_128246560, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128246112_128246336, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer4_128123904_128124128);
   U1210 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263672_128263840);
   U1211 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263672_128263840);
   U1212 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263672_128263840);
   U1213 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263672_128263840);
   U1214 : XOR2X1 port map( A => n3923, B => n917, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_11_port);
   U1215 : XOR2X1 port map( A => n3966, B => n1076, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_11_port);
   U1216 : XOR2X1 port map( A => n4052, B => n599, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_11_port);
   U1217 : XOR2X1 port map( A => n3880, B => n758, Y => 
                           input_times_b0_div_componentxinput_A_inverted_11_port);
   U1218 : XOR2X1 port map( A => n3922, B => n899, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_13_port);
   U1219 : XOR2X1 port map( A => n3965, B => n1058, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_13_port);
   U1220 : XOR2X1 port map( A => n4051, B => n581, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_13_port);
   U1221 : XOR2X1 port map( A => n3879, B => n740, Y => 
                           input_times_b0_div_componentxinput_A_inverted_13_port);
   U1222 : XNOR2X1 port map( A => n43, B => n908, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_12_port);
   U1223 : NOR2X1 port map( A => n3923, B => n917, Y => n43);
   U1224 : XNOR2X1 port map( A => n44, B => n1067, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_12_port);
   U1225 : NOR2X1 port map( A => n3966, B => n1076, Y => n44);
   U1226 : XNOR2X1 port map( A => n45, B => n590, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_12_port);
   U1227 : NOR2X1 port map( A => n4052, B => n599, Y => n45);
   U1228 : XNOR2X1 port map( A => n46, B => n749, Y => 
                           input_times_b0_div_componentxinput_A_inverted_12_port);
   U1229 : NOR2X1 port map( A => n3880, B => n758, Y => n46);
   U1230 : XOR2X1 port map( A => n3924, B => n930, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_10_port);
   U1231 : NAND2X1 port map( A => n3914, B => n4441, Y => n3924);
   U1232 : XOR2X1 port map( A => n3967, B => n1089, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_10_port);
   U1233 : NAND2X1 port map( A => n3957, B => n4494, Y => n3967);
   U1234 : XOR2X1 port map( A => n4053, B => n612, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_10_port);
   U1235 : NAND2X1 port map( A => n4043, B => n4600, Y => n4053);
   U1236 : XOR2X1 port map( A => n3881, B => n771, Y => 
                           input_times_b0_div_componentxinput_A_inverted_10_port);
   U1237 : NAND2X1 port map( A => n3871, B => input_times_b0_mul_componentxn90,
                           Y => n3881);
   U1238 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128263672_128263840, B 
                           => n2835, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128237752_128237976_128238144);
   U1239 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128263672_128263840);
   U1240 : XOR2X1 port map( A => n880, B => n878, Y => n2835);
   U1241 : INVX1 port map( A => n2810, Y => n880);
   U1242 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128263672_128263840, B 
                           => n3069, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128237752_128237976_128238144);
   U1243 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128263672_128263840);
   U1244 : XOR2X1 port map( A => n1039, B => n1037, Y => n3069);
   U1245 : INVX1 port map( A => n3044, Y => n1039);
   U1246 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128263672_128263840, B 
                           => n3537, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128237752_128237976_128238144);
   U1247 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128263672_128263840);
   U1248 : XOR2X1 port map( A => n562, B => n560, Y => n3537);
   U1249 : INVX1 port map( A => n3512, Y => n562);
   U1250 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128263672_128263840, B 
                           => n2601, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128237752_128237976_128238144);
   U1251 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198976_128199144, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198472_128198640_128198808, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128263672_128263840);
   U1252 : XOR2X1 port map( A => n721, B => n719, Y => n2601);
   U1253 : INVX1 port map( A => n2576, Y => n721);
   U1254 : INVX1 port map( A => n2812, Y => n878);
   U1255 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_128198024_128197968, 
                           B0 => n2811, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198080_128198192_128198360, Y 
                           => n2812);
   U1256 : INVX1 port map( A => n3046, Y => n1037);
   U1257 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_128198024_128197968, 
                           B0 => n3045, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198080_128198192_128198360, Y 
                           => n3046);
   U1258 : INVX1 port map( A => n3514, Y => n560);
   U1259 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_128198024_128197968, 
                           B0 => n3513, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198080_128198192_128198360, Y 
                           => n3514);
   U1260 : INVX1 port map( A => n2578, Y => n719);
   U1261 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197464_128197688_128197856, 
                           A1 => 
                           input_times_b0_mul_componentxUMxcarry_layer2_128198024_128197968, 
                           B0 => n2577, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198080_128198192_128198360, Y 
                           => n2578);
   U1262 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_3_port);
   U1263 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_3_port);
   U1264 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_3_port);
   U1265 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127672448_127826240_127826520, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127826128_127826296, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_3_port)
                           ;
   U1266 : OR3XL port map( A => n986, B => n980, C => n3917, Y => n3916);
   U1267 : OR3XL port map( A => n1145, B => n1139, C => n3960, Y => n3959);
   U1268 : OR3XL port map( A => n668, B => n662, C => n4046, Y => n4045);
   U1269 : OR3XL port map( A => n827, B => n821, C => n3874, Y => n3873);
   U1270 : INVX1 port map( A => n4441, Y => n940);
   U1271 : INVX1 port map( A => n4494, Y => n1099);
   U1272 : INVX1 port map( A => n4600, Y => n622);
   U1273 : INVX1 port map( A => input_times_b0_mul_componentxn90, Y => n781);
   U1274 : XOR2X1 port map( A => n3915, B => n957, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_7_port);
   U1275 : XOR2X1 port map( A => n3958, B => n1116, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_7_port);
   U1276 : XOR2X1 port map( A => n4044, B => n639, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_7_port);
   U1277 : XOR2X1 port map( A => n3872, B => n798, Y => 
                           input_times_b0_div_componentxinput_A_inverted_7_port
                           );
   U1278 : XNOR2X1 port map( A => n47, B => n950, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_8_port);
   U1279 : NOR2X1 port map( A => n957, B => n3915, Y => n47);
   U1280 : XNOR2X1 port map( A => n48, B => n1109, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_8_port);
   U1281 : NOR2X1 port map( A => n1116, B => n3958, Y => n48);
   U1282 : XNOR2X1 port map( A => n49, B => n632, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_8_port);
   U1283 : NOR2X1 port map( A => n639, B => n4044, Y => n49);
   U1284 : XNOR2X1 port map( A => n50, B => n791, Y => 
                           input_times_b0_div_componentxinput_A_inverted_8_port
                           );
   U1285 : NOR2X1 port map( A => n798, B => n3872, Y => n50);
   U1286 : XOR2X1 port map( A => n3916, B => n972, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_5_port);
   U1287 : XOR2X1 port map( A => n3959, B => n1131, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_5_port);
   U1288 : XOR2X1 port map( A => n4045, B => n654, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_5_port);
   U1289 : XOR2X1 port map( A => n3873, B => n813, Y => 
                           input_times_b0_div_componentxinput_A_inverted_5_port
                           );
   U1290 : XNOR2X1 port map( A => n51, B => n965, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_6_port);
   U1291 : NOR2X1 port map( A => n972, B => n3916, Y => n51);
   U1292 : XNOR2X1 port map( A => n52, B => n1124, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_6_port);
   U1293 : NOR2X1 port map( A => n1131, B => n3959, Y => n52);
   U1294 : XNOR2X1 port map( A => n53, B => n647, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_6_port);
   U1295 : NOR2X1 port map( A => n654, B => n4045, Y => n53);
   U1296 : XNOR2X1 port map( A => n54, B => n806, Y => 
                           input_times_b0_div_componentxinput_A_inverted_6_port
                           );
   U1297 : NOR2X1 port map( A => n813, B => n3873, Y => n54);
   U1298 : BUFX3 port map( A => n81, Y => n126);
   U1299 : BUFX3 port map( A => n82, Y => n130);
   U1300 : BUFX3 port map( A => n83, Y => n118);
   U1301 : BUFX3 port map( A => n84, Y => n122);
   U1302 : BUFX3 port map( A => n81, Y => n125);
   U1303 : BUFX3 port map( A => n82, Y => n129);
   U1304 : BUFX3 port map( A => n83, Y => n117);
   U1305 : BUFX3 port map( A => n84, Y => n121);
   U1306 : XOR2X1 port map( A => n3917, B => n986, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_3_port);
   U1307 : XOR2X1 port map( A => n3960, B => n1145, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_3_port);
   U1308 : XOR2X1 port map( A => n4046, B => n668, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_3_port);
   U1309 : XOR2X1 port map( A => n3874, B => n827, Y => 
                           input_times_b0_div_componentxinput_A_inverted_3_port
                           );
   U1310 : XNOR2X1 port map( A => n55, B => n980, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_4_port);
   U1311 : NOR2X1 port map( A => n986, B => n3917, Y => n55);
   U1312 : XNOR2X1 port map( A => n56, B => n1139, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_4_port);
   U1313 : NOR2X1 port map( A => n1145, B => n3960, Y => n56);
   U1314 : XNOR2X1 port map( A => n57, B => n662, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_4_port);
   U1315 : NOR2X1 port map( A => n668, B => n4046, Y => n57);
   U1316 : XNOR2X1 port map( A => n58, B => n821, Y => 
                           input_times_b0_div_componentxinput_A_inverted_4_port
                           );
   U1317 : NOR2X1 port map( A => n827, B => n3874, Y => n58);
   U1318 : NAND3BX1 port map( AN => output_contracterxn6, B => 
                           output_previous_1_8_port, C => 
                           output_previous_1_9_port, Y => output_contracterxn3)
                           ;
   U1319 : NAND3BX1 port map( AN => output_contracterxn5, B => 
                           output_previous_1_13_port, C => 
                           output_previous_1_14_port, Y => output_contracterxn4
                           );
   U1320 : NOR3X1 port map( A => output_contracterxn8, B => 
                           output_previous_1_11_port, C => 
                           output_previous_1_10_port, Y => output_contracterxn1
                           );
   U1321 : NOR3X1 port map( A => results_a1_a2_7_port, B => 
                           results_a1_a2_8_port, C => 
                           results_a1_a2_inv_inverterxn4, Y => 
                           results_a1_a2_inv_inverterxn2);
   U1322 : AOI22X1 port map( A0 => results_a1_a2_inv_3_port, A1 => 
                           results_b0_b1_b2_3_port, B0 => n4164, B1 => n4165, Y
                           => n4163);
   U1323 : AOI22X1 port map( A0 => results_a1_a2_inv_5_port, A1 => 
                           results_b0_b1_b2_5_port, B0 => n4160, B1 => n4161, Y
                           => n4159);
   U1324 : AOI22X1 port map( A0 => results_a1_a2_inv_7_port, A1 => 
                           results_b0_b1_b2_7_port, B0 => n4156, B1 => n4157, Y
                           => n4155);
   U1325 : AOI22X1 port map( A0 => results_a1_a2_inv_9_port, A1 => 
                           results_b0_b1_b2_9_port, B0 => n4152, B1 => n4153, Y
                           => n4183);
   U1326 : AOI22X1 port map( A0 => results_a1_a2_inv_11_port, A1 => 
                           results_b0_b1_b2_11_port, B0 => n4181, B1 => n4182, 
                           Y => n4179);
   U1327 : AOI22X1 port map( A0 => results_a1_a2_inv_13_port, A1 => 
                           results_b0_b1_b2_13_port, B0 => n4177, B1 => n4178, 
                           Y => n4175);
   U1328 : OAI2BB2X1 port map( B0 => n4167, B1 => n4166, A0N => 
                           results_a1_a2_inv_2_port, A1N => 
                           results_b0_b1_b2_2_port, Y => n4164);
   U1329 : OAI2BB2X1 port map( B0 => n4163, B1 => n4162, A0N => 
                           results_a1_a2_inv_4_port, A1N => 
                           results_b0_b1_b2_4_port, Y => n4160);
   U1330 : OAI2BB2X1 port map( B0 => n4159, B1 => n4158, A0N => 
                           results_a1_a2_inv_6_port, A1N => 
                           results_b0_b1_b2_6_port, Y => n4156);
   U1331 : OAI2BB2X1 port map( B0 => n4155, B1 => n4154, A0N => 
                           results_a1_a2_inv_8_port, A1N => 
                           results_b0_b1_b2_8_port, Y => n4152);
   U1332 : OAI2BB2X1 port map( B0 => n4183, B1 => n4184, A0N => 
                           results_a1_a2_inv_10_port, A1N => 
                           results_b0_b1_b2_10_port, Y => n4181);
   U1333 : OAI2BB2X1 port map( B0 => n4179, B1 => n4180, A0N => 
                           results_a1_a2_inv_12_port, A1N => 
                           results_b0_b1_b2_12_port, Y => n4177);
   U1334 : OAI2BB2X1 port map( B0 => n4175, B1 => n4176, A0N => 
                           results_a1_a2_inv_14_port, A1N => 
                           results_b0_b1_b2_14_port, Y => n4173);
   U1335 : INVX1 port map( A => n3192, Y => n497);
   U1336 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127672560_127674464, 
                           A1 => n501, B0 => n3191, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830672_127844928_127846832, Y 
                           => n3192);
   U1337 : XNOR2X1 port map( A => results_a1_a2_inv_inverterxn2, B => 
                           results_a1_a2_9_port, Y => results_a1_a2_inv_9_port)
                           ;
   U1338 : XOR2X1 port map( A => n513, B => n3193, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127731808_127826912_127827136);
   U1339 : XOR2X1 port map( A => results_b0_b1_b2_3_port, B => 
                           results_a1_a2_inv_3_port, Y => n4165);
   U1340 : XOR2X1 port map( A => results_b0_b1_b2_5_port, B => 
                           results_a1_a2_inv_5_port, Y => n4161);
   U1341 : XOR2X1 port map( A => results_b0_b1_b2_7_port, B => 
                           results_a1_a2_inv_7_port, Y => n4157);
   U1342 : XOR2X1 port map( A => results_b0_b1_b2_9_port, B => 
                           results_a1_a2_inv_9_port, Y => n4153);
   U1343 : XOR2X1 port map( A => results_b0_b1_b2_11_port, B => 
                           results_a1_a2_inv_11_port, Y => n4182);
   U1344 : XOR2X1 port map( A => results_b0_b1_b2_13_port, B => 
                           results_a1_a2_inv_13_port, Y => n4178);
   U1345 : XOR2X1 port map( A => results_b0_b1_b2_15_port, B => 
                           results_a1_a2_inv_15_port, Y => n4174);
   U1346 : XOR2X1 port map( A => n501, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127672560_127674464, Y 
                           => n3191);
   U1347 : XOR2X1 port map( A => n493, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127827304_127827416, Y 
                           => n3251);
   U1348 : OR3XL port map( A => results_a1_a2_5_port, B => results_a1_a2_6_port
                           , C => results_a1_a2_inv_inverterxn6, Y => 
                           results_a1_a2_inv_inverterxn4);
   U1349 : BUFX3 port map( A => n4557, Y => n232);
   U1350 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_17,
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_17_port, 
                           B1 => n4548, Y => n4557);
   U1351 : XOR2X1 port map( A => n3815, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_17,
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_17_port);
   U1352 : XOR2X1 port map( A => n2354, B => n2355, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_17)
                           ;
   U1353 : XNOR2X1 port map( A => results_b0_b1_b2_2_port, B => 
                           results_a1_a2_inv_2_port, Y => n4166);
   U1354 : XNOR2X1 port map( A => results_b0_b1_b2_4_port, B => 
                           results_a1_a2_inv_4_port, Y => n4162);
   U1355 : XNOR2X1 port map( A => results_b0_b1_b2_6_port, B => 
                           results_a1_a2_inv_6_port, Y => n4158);
   U1356 : XNOR2X1 port map( A => results_b0_b1_b2_8_port, B => 
                           results_a1_a2_inv_8_port, Y => n4154);
   U1357 : XNOR2X1 port map( A => results_b0_b1_b2_10_port, B => 
                           results_a1_a2_inv_10_port, Y => n4184);
   U1358 : XNOR2X1 port map( A => results_b0_b1_b2_12_port, B => 
                           results_a1_a2_inv_12_port, Y => n4180);
   U1359 : XNOR2X1 port map( A => results_b0_b1_b2_14_port, B => 
                           results_a1_a2_inv_14_port, Y => n4176);
   U1360 : BUFX3 port map( A => n4546, Y => n231);
   U1361 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_0_port, 
                           A1 => n133, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_0_port, 
                           B1 => n165, Y => n4546);
   U1362 : BUFX3 port map( A => n4538, Y => n230);
   U1363 : AOI22XL port map( A0 => output_signal_1_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_1_port, 
                           B1 => n165, Y => n4538);
   U1364 : XOR2X1 port map( A => output_signal_1_port, B => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_0_port, Y 
                           => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_1_port);
   U1365 : INVX1 port map( A => n165, Y => n1203);
   U1366 : INVX1 port map( A => n4172, Y => n1205);
   U1367 : AOI22X1 port map( A0 => results_a1_a2_inv_15_port, A1 => 
                           results_b0_b1_b2_15_port, B0 => n4173, B1 => n4174, 
                           Y => n4172);
   U1368 : INVX1 port map( A => n3252, Y => n482);
   U1369 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127827304_127827416, 
                           A1 => n493, B0 => n3251, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827248_127827472_127827640, Y 
                           => n3252);
   U1370 : AOI22X1 port map( A0 => output_previous_1_10_port, A1 => n133, B0 =>
                           output_p1_times_a1_mul_componentxinput_A_inverted_10_port, 
                           B1 => n165, Y => n4545);
   U1371 : XOR2X1 port map( A => n3790, B => output_previous_1_10_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_10_port);
   U1372 : NAND2X1 port map( A => n3775, B => n1210, Y => n3790);
   U1373 : AOI22X1 port map( A0 => output_previous_1_11_port, A1 => n133, B0 =>
                           output_p1_times_a1_mul_componentxinput_A_inverted_11_port, 
                           B1 => n165, Y => n4544);
   U1374 : XOR2X1 port map( A => n3788, B => output_previous_1_11_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_11_port);
   U1375 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_9, 
                           A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_9_port, 
                           B1 => n4548, Y => n4547);
   U1376 : XNOR2X1 port map( A => n3807, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_9, 
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_9_port);
   U1377 : NOR3X1 port map( A => results_a1_a2_13_port, B => 
                           results_a1_a2_14_port, C => 
                           results_a1_a2_inv_inverterxn13, Y => 
                           results_a1_a2_inv_inverterxn12);
   U1378 : INVX1 port map( A => n3122, Y => n450);
   U1379 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b9, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b10, B0 
                           => n3121, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b8, Y => 
                           n3122);
   U1380 : INVX1 port map( A => n4561, Y => n423);
   U1381 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_13,
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_13_port, 
                           B1 => n4548, Y => n4561);
   U1382 : XOR2X1 port map( A => n3818, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_13,
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_13_port);
   U1383 : INVX1 port map( A => n4558, Y => n401);
   U1384 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_16,
                           A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_16_port, 
                           B1 => n4548, Y => n4558);
   U1385 : XNOR2X1 port map( A => n3816, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_16,
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_16_port);
   U1386 : INVX1 port map( A => n3204, Y => n461);
   U1387 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
                           A1 => n512, B0 => n3203, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673120_127675024_127730240, Y 
                           => n3204);
   U1388 : INVX1 port map( A => n3216, Y => n434);
   U1389 : AOI22X1 port map( A0 => n511, A1 => n491, B0 => n3215, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831456_127845712_127847616, Y 
                           => n3216);
   U1390 : INVX1 port map( A => n3218, Y => n456);
   U1391 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
                           B0 => n3217, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635920_127637824_127713520, Y 
                           => n3218);
   U1392 : INVX1 port map( A => n3116, Y => n458);
   U1393 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b8, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b9, B0 =>
                           n3115, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b7, Y => 
                           n3116);
   U1394 : INVX1 port map( A => n3206, Y => n457);
   U1395 : AOI22X1 port map( A0 => n486, A1 => n458, B0 => n3205, B1 => n505, Y
                           => n3206);
   U1396 : NAND3BX1 port map( AN => results_a1_a2_10_port, B => n1302, C => 
                           results_a1_a2_inv_inverterxn2, Y => 
                           results_a1_a2_inv_inverterxn15);
   U1397 : NOR2BX1 port map( AN => results_a1_a2_inv_inverterxn12, B => 
                           results_a1_a2_15_port, Y => 
                           results_a1_a2_inv_inverterxn11);
   U1398 : XNOR2X1 port map( A => results_a1_a2_inv_inverterxn12, B => 
                           results_a1_a2_15_port, Y => 
                           results_a1_a2_inv_15_port);
   U1399 : XNOR2X1 port map( A => results_a1_a2_inv_inverterxn11, B => 
                           results_a1_a2_16_port, Y => 
                           results_a1_a2_inv_16_port);
   U1400 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b11
                           , B => n3143, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831568_127845824_127847728);
   U1401 : XOR2X1 port map( A => results_a1_a2_inv_inverterxn15, B => 
                           results_a1_a2_11_port, Y => 
                           results_a1_a2_inv_11_port);
   U1402 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b7,
                           B => n3115, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831120_127845376_127847280);
   U1403 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b9,
                           B => n3127, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831344_127845600_127847504);
   U1404 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b10
                           , B => output_p1_times_a1_mul_componentxUMxa1_and_b9
                           , Y => n3121);
   U1405 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b11
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b10, Y =>
                           n3127);
   U1406 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b12
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b11, Y =>
                           n3135);
   U1407 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b13
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b12, Y =>
                           n3143);
   U1408 : XOR2X1 port map( A => results_a1_a2_inv_inverterxn13, B => 
                           results_a1_a2_13_port, Y => 
                           results_a1_a2_inv_13_port);
   U1409 : XOR2X1 port map( A => results_a1_a2_inv_inverterxn4, B => 
                           results_a1_a2_7_port, Y => results_a1_a2_inv_7_port)
                           ;
   U1410 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b8,
                           B => output_p1_times_a1_mul_componentxUMxa1_and_b7, 
                           Y => n3109);
   U1411 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b9,
                           B => output_p1_times_a1_mul_componentxUMxa1_and_b8, 
                           Y => n3115);
   U1412 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b9,
                           B => output_p1_times_a1_mul_componentxUMxa4_and_b8, 
                           Y => n3137);
   U1413 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b8,
                           B => output_p1_times_a1_mul_componentxUMxa4_and_b7, 
                           Y => n3129);
   U1414 : XOR2X1 port map( A => results_a1_a2_inv_inverterxn8, B => 
                           results_a1_a2_3_port, Y => results_a1_a2_inv_3_port)
                           ;
   U1415 : XOR2X1 port map( A => results_a1_a2_inv_inverterxn6, B => 
                           results_a1_a2_5_port, Y => results_a1_a2_inv_5_port)
                           ;
   U1416 : XOR2X1 port map( A => n508, B => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830560_127844816_127846720, Y 
                           => n3189);
   U1417 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831008_127845264_127847168, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673008_127674912_127730128, Y 
                           => n3199);
   U1418 : XOR2X1 port map( A => n512, B => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831120_127845376_127847280, Y 
                           => n3203);
   U1419 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831232_127845488_127847392, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673232_127675136_127730352, Y 
                           => n3207);
   U1420 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673456_127675360_127730576, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732480_127722160_127724064, Y 
                           => n3217);
   U1421 : XOR2X1 port map( A => n504, B => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831568_127845824_127847728, Y 
                           => n3221);
   U1422 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127635696_127637600, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831344_127845600_127847504, Y 
                           => n3211);
   U1423 : XOR2X1 port map( A => n479, B => n500, Y => n3197);
   U1424 : XOR2X1 port map( A => n487, B => n506, Y => n3195);
   U1425 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672672_127674576_127729792, B 
                           => n502, Y => n3247);
   U1426 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732144_127721824_127723728, B 
                           => n477, Y => n3255);
   U1427 : XOR2X1 port map( A => n491, B => n511, Y => n3215);
   U1428 : XOR2X1 port map( A => n458, B => n486, Y => n3205);
   U1429 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635696_127637600, B 
                           => n468, Y => n3257);
   U1430 : XOR2X1 port map( A => n450, B => n476, Y => n3209);
   U1431 : XOR2X1 port map( A => n435, B => n434, Y => n3265);
   U1432 : OR3XL port map( A => results_a1_a2_11_port, B => 
                           results_a1_a2_12_port, C => 
                           results_a1_a2_inv_inverterxn15, Y => 
                           results_a1_a2_inv_inverterxn13);
   U1433 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127827304_127827416);
   U1434 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127827752_127827920);
   U1435 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b8,
                           B => n3121, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831232_127845488_127847392);
   U1436 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b7,
                           B => n3137, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673456_127675360_127730576);
   U1437 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827752_127827920);
   U1438 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732032_127721712_127723616, B 
                           => n3199, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221424_128221536_128221704);
   U1439 : XOR2X1 port map( A => n467, B => n3213, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127715424_128223048_128223272);
   U1440 : XNOR2X1 port map( A => n59, B => results_a1_a2_4_port, Y => 
                           results_a1_a2_inv_4_port);
   U1441 : NOR2X1 port map( A => results_a1_a2_3_port, B => 
                           results_a1_a2_inv_inverterxn8, Y => n59);
   U1442 : XNOR2X1 port map( A => n60, B => results_a1_a2_6_port, Y => 
                           results_a1_a2_inv_6_port);
   U1443 : NOR2X1 port map( A => results_a1_a2_5_port, B => 
                           results_a1_a2_inv_inverterxn6, Y => n60);
   U1444 : XNOR2X1 port map( A => n61, B => results_a1_a2_8_port, Y => 
                           results_a1_a2_inv_8_port);
   U1445 : NOR2X1 port map( A => results_a1_a2_7_port, B => 
                           results_a1_a2_inv_inverterxn4, Y => n61);
   U1446 : XOR2X1 port map( A => results_a1_a2_inv_inverterxn17, B => 
                           results_a1_a2_10_port, Y => 
                           results_a1_a2_inv_10_port);
   U1447 : NAND2X1 port map( A => results_a1_a2_inv_inverterxn2, B => n1302, Y 
                           => results_a1_a2_inv_inverterxn17);
   U1448 : XNOR2X1 port map( A => n62, B => results_a1_a2_12_port, Y => 
                           results_a1_a2_inv_12_port);
   U1449 : NOR2X1 port map( A => results_a1_a2_inv_inverterxn15, B => 
                           results_a1_a2_11_port, Y => n62);
   U1450 : XNOR2X1 port map( A => n63, B => results_a1_a2_14_port, Y => 
                           results_a1_a2_inv_14_port);
   U1451 : NOR2X1 port map( A => results_a1_a2_13_port, B => 
                           results_a1_a2_inv_inverterxn13, Y => n63);
   U1452 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b10
                           , B => n3135, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831456_127845712_127847616);
   U1453 : XOR2X1 port map( A => results_b0_b1_b2_16_port, B => 
                           results_a1_a2_inv_16_port, Y => n4171);
   U1454 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827304_127827416);
   U1455 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830896_127845152_127847056, B 
                           => n3195, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827248_127827472_127827640);
   U1456 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830672_127844928_127846832, B 
                           => n3191, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127826576_127826800_127826968);
   U1457 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127731920_127721600, B 
                           => n3197, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127827584_127827808_128221256);
   U1458 : XOR2X1 port map( A => n499, B => n3209, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222376_128222600_128222768);
   U1459 : OR3XL port map( A => results_a1_a2_3_port, B => results_a1_a2_4_port
                           , C => results_a1_a2_inv_inverterxn8, Y => 
                           results_a1_a2_inv_inverterxn6);
   U1460 : XOR2X1 port map( A => n492, B => n3201, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127635584_128221368_128221592);
   U1461 : XOR2X1 port map( A => n505, B => n3205, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221872_128222096_128222264);
   U1462 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673344_127675248_127730464, B 
                           => n3211, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222936_128223104_128223216);
   U1463 : INVX1 port map( A => n4550, Y => n480);
   U1464 : AOI22X1 port map( A0 => n2353, A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_7_port, 
                           B1 => n4548, Y => n4550);
   U1465 : XOR2X1 port map( A => n3809, B => n2353, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_7_port);
   U1466 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n510, Y => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer3_128246112_128246336);
   U1467 : BUFX3 port map( A => n4537, Y => n229);
   U1468 : AOI22X1 port map( A0 => output_signal_2_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_2_port, 
                           B1 => n165, Y => n4537);
   U1469 : XNOR2X1 port map( A => output_signal_2_port, B => n3782, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_2_port);
   U1470 : NOR2XL port map( A => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_0_port, B 
                           => output_signal_1_port, Y => n3782);
   U1471 : INVX1 port map( A => n4559, Y => n408);
   U1472 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_15,
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_15_port, 
                           B1 => n4548, Y => n4559);
   U1473 : XNOR2X1 port map( A => n3817, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_15,
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_15_port);
   U1474 : INVX1 port map( A => n4549, Y => n473);
   U1475 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_8, 
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_8_port, 
                           B1 => n4548, Y => n4549);
   U1476 : XOR2X1 port map( A => n3808, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_8, 
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_8_port);
   U1477 : OR2X2 port map( A => n2353, B => n3809, Y => n3808);
   U1478 : INVX1 port map( A => n4560, Y => n417);
   U1479 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_14,
                           A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_14_port, 
                           B1 => n4548, Y => n4560);
   U1480 : XOR2X1 port map( A => n3819, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_14,
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_14_port);
   U1481 : OR2X2 port map( A => 
                           output_p1_times_a1_mul_componentxunsigned_output_13,
                           B => n3818, Y => n3819);
   U1482 : BUFX3 port map( A => n4536, Y => n228);
   U1483 : AOI22X1 port map( A0 => output_signal_3_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_3_port, 
                           B1 => n165, Y => n4536);
   U1484 : XOR2X1 port map( A => n3781, B => output_signal_3_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_3_port);
   U1485 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672560_127674464, B 
                           => n3189, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127826464_127826632_127826744);
   U1486 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830448_127844704_127846608, B 
                           => n3187, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127672448_127826240_127826520);
   U1487 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673120_127675024_127730240, B 
                           => n3203, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128221760_128221928_128222040);
   U1488 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732256_127721936_127723840, B 
                           => n3207, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128222432_128222544_128222712);
   U1489 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n510, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128246112_128246336);
   U1490 : BUFX3 port map( A => n4535, Y => n227);
   U1491 : AOI22X1 port map( A0 => output_signal_4_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_4_port, 
                           B1 => n165, Y => n4535);
   U1492 : XOR2X1 port map( A => n3780, B => output_signal_4_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_4_port);
   U1493 : OR2X2 port map( A => output_signal_3_port, B => n3781, Y => n3780);
   U1494 : INVX1 port map( A => n4562, Y => n432);
   U1495 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_12,
                           A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_12_port, 
                           B1 => n4548, Y => n4562);
   U1496 : XOR2X1 port map( A => n3821, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_12,
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_12_port);
   U1497 : OR2X2 port map( A => n3820, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_11,
                           Y => n3821);
   U1498 : INVX1 port map( A => n4564, Y => n453);
   U1499 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_10,
                           A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_10_port, 
                           B1 => n4548, Y => n4564);
   U1500 : XOR2X1 port map( A => n3822, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_10,
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_10_port);
   U1501 : NAND2X1 port map( A => n3807, B => n462, Y => n3822);
   U1502 : BUFX3 port map( A => n4534, Y => n226);
   U1503 : AOI22X1 port map( A0 => output_signal_5_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_5_port, 
                           B1 => n165, Y => n4534);
   U1504 : XOR2X1 port map( A => n3779, B => output_signal_5_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_5_port);
   U1505 : BUFX3 port map( A => n4533, Y => n225);
   U1506 : AOI22X1 port map( A0 => output_signal_6_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_6_port, 
                           B1 => n165, Y => n4533);
   U1507 : XOR2X1 port map( A => n3778, B => output_signal_6_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_6_port);
   U1508 : OR2X2 port map( A => output_signal_5_port, B => n3779, Y => n3778);
   U1509 : INVX1 port map( A => n3128, Y => n436);
   U1510 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b10, A1 
                           => output_p1_times_a1_mul_componentxUMxa0_and_b11, 
                           B0 => n3127, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b9, Y => 
                           n3128);
   U1511 : INVX1 port map( A => n3190, Y => n502);
   U1512 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
                           A1 => n508, B0 => n3189, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672560_127674464, Y 
                           => n3190);
   U1513 : INVX1 port map( A => n3198, Y => n477);
   U1514 : AOI22X1 port map( A0 => n500, A1 => n479, B0 => n3197, B1 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127731920_127721600, Y 
                           => n3198);
   U1515 : INVX1 port map( A => n3208, Y => n451);
   U1516 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
                           B0 => n3207, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732256_127721936_127723840, Y 
                           => n3208);
   U1517 : INVX1 port map( A => n3212, Y => n439);
   U1518 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127635696_127637600, 
                           B0 => n3211, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673344_127675248_127730464, Y 
                           => n3212);
   U1519 : INVX1 port map( A => n3266, Y => n433);
   U1520 : AOI22X1 port map( A0 => n434, A1 => n435, B0 => n3265, B1 => n456, Y
                           => n3266);
   U1521 : BUFX3 port map( A => n4532, Y => n224);
   U1522 : AOI22X1 port map( A0 => output_signal_7_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_7_port, 
                           B1 => n165, Y => n4532);
   U1523 : XOR2X1 port map( A => n3777, B => output_signal_7_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_7_port);
   U1524 : INVX1 port map( A => n4563, Y => n441);
   U1525 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_11,
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_11_port, 
                           B1 => n4548, Y => n4563);
   U1526 : XOR2X1 port map( A => n3820, B => 
                           output_p1_times_a1_mul_componentxunsigned_output_11,
                           Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_11_port);
   U1527 : INVX1 port map( A => n3196, Y => n483);
   U1528 : AOI22X1 port map( A0 => n506, A1 => n487, B0 => n3195, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830896_127845152_127847056, Y 
                           => n3196);
   U1529 : INVX1 port map( A => n3256, Y => n470);
   U1530 : AOI22X1 port map( A0 => n477, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
                           B0 => n3255, B1 => n471, Y => n3256);
   U1531 : INVX1 port map( A => n3258, Y => n459);
   U1532 : AOI22X1 port map( A0 => n468, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635696_127637600, 
                           B0 => n3257, B1 => n461, Y => n3258);
   U1533 : INVX1 port map( A => n3210, Y => n447);
   U1534 : AOI22X1 port map( A0 => n476, A1 => n450, B0 => n3209, B1 => n499, Y
                           => n3210);
   U1535 : BUFX3 port map( A => n4531, Y => n223);
   U1536 : AOI22X1 port map( A0 => output_previous_1_8_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_8_port, 
                           B1 => n165, Y => n4531);
   U1537 : XOR2X1 port map( A => n3776, B => output_previous_1_8_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_8_port);
   U1538 : OR2X2 port map( A => output_signal_7_port, B => n3777, Y => n3776);
   U1539 : INVX1 port map( A => n3200, Y => n471);
   U1540 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
                           B0 => n3199, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732032_127721712_127723616, Y 
                           => n3200);
   U1541 : INVX1 port map( A => n3248, Y => n496);
   U1542 : AOI22X1 port map( A0 => n502, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
                           B0 => n3247, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127826576_127826800_127826968, Y 
                           => n3248);
   U1543 : BUFX3 port map( A => n4530, Y => n222);
   U1544 : AOI22X1 port map( A0 => output_previous_1_9_port, A1 => n134, B0 => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_9_port, 
                           B1 => n165, Y => n4530);
   U1545 : XNOR2X1 port map( A => n3775, B => output_previous_1_9_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_9_port);
   U1546 : INVX1 port map( A => results_a1_a2_9_port, Y => n1302);
   U1547 : AOI22X1 port map( A0 => output_previous_1_12_port, A1 => n133, B0 =>
                           output_p1_times_a1_mul_componentxinput_A_inverted_12_port, 
                           B1 => n165, Y => n4543);
   U1548 : XOR2X1 port map( A => n3789, B => output_previous_1_12_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_12_port);
   U1549 : OR2X2 port map( A => n3788, B => output_previous_1_11_port, Y => 
                           n3789);
   U1550 : AOI22X1 port map( A0 => output_previous_1_13_port, A1 => n133, B0 =>
                           output_p1_times_a1_mul_componentxinput_A_inverted_13_port, 
                           B1 => n165, Y => n4542);
   U1551 : XOR2X1 port map( A => n3786, B => output_previous_1_13_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_13_port);
   U1552 : INVX1 port map( A => n3136, Y => n428);
   U1553 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b11, A1 
                           => output_p1_times_a1_mul_componentxUMxa0_and_b12, 
                           B0 => n3135, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b10, Y =>
                           n3136);
   U1554 : INVX1 port map( A => n3146, Y => n446);
   U1555 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b9, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b10, B0 
                           => n3145, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b8, Y => 
                           n3146);
   U1556 : INVX1 port map( A => n3144, Y => n426);
   U1557 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b12, A1 
                           => output_p1_times_a1_mul_componentxUMxa0_and_b13, 
                           B0 => n3143, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b11, Y =>
                           n3144);
   U1558 : INVX1 port map( A => n4552, Y => n495);
   U1559 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_5_port, 
                           A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_5_port, 
                           B1 => n4548, Y => n4552);
   U1560 : XOR2X1 port map( A => n3811, B => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_5_port, Y 
                           => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_5_port);
   U1561 : INVX1 port map( A => n3228, Y => n442);
   U1562 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127715536_127848576, 
                           A1 => n498, B0 => n3227, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831680_127845936_127847840, Y 
                           => n3228);
   U1563 : AOI22X1 port map( A0 => n507, A1 => n484, B0 => n3239, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831904_127846160_127848064, Y 
                           => n3240);
   U1564 : INVX1 port map( A => n3138, Y => n455);
   U1565 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b8, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b9, B0 =>
                           n3137, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b7, Y => 
                           n3138);
   U1566 : INVX1 port map( A => n3234, Y => n465);
   U1567 : AOI22X1 port map( A0 => n490, A1 => n466, B0 => n3233, B1 => n514, Y
                           => n3234);
   U1568 : OR3XL port map( A => output_signal_1_port, B => output_signal_2_port
                           , C => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_0_port, Y 
                           => n3781);
   U1569 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_2_port);
   U1570 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b10
                           , B => n3163, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673792_127675696_127730912);
   U1571 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b10
                           , B => output_p1_times_a1_mul_componentxUMxa4_and_b9
                           , Y => n3145);
   U1572 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b11
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b10, Y =>
                           n3153);
   U1573 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b12
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b11, Y =>
                           n3163);
   U1574 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b14
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b13, Y =>
                           n3151);
   U1575 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b15
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b14, Y =>
                           n3161);
   U1576 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b8,
                           B => output_p1_times_a1_mul_componentxUMxa7_and_b7, 
                           Y => n3155);
   U1577 : XOR2X1 port map( A => n474, B => n3225, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224392_128224616_128224784);
   U1578 : XOR2X1 port map( A => n514, B => n3233, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128197016_128197240_128197352);
   U1579 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732592_127722272_127724176, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636032_127637936_127713632, Y 
                           => n3223);
   U1580 : XOR2X1 port map( A => n498, B => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127715536_127848576, Y 
                           => n3227);
   U1581 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673680_127675584_127730800, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732704_127722384_127724288, Y 
                           => n3229);
   U1582 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715648_127848688_127850592, B 
                           => n427, Y => n3269);
   U1583 : XOR2X1 port map( A => n466, B => n490, Y => n3233);
   U1584 : XOR2X1 port map( A => n484, B => n507, Y => n3239);
   U1585 : XOR2X1 port map( A => n410, B => n465, Y => n3277);
   U1586 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b13
                           , B => n3161, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831792_127846048_127847952);
   U1587 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b9,
                           B => n3153, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673680_127675584_127730800);
   U1588 : XOR2X1 port map( A => n485, B => n3219, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223720_128223944_128224168);
   U1589 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636144_127638048_127713744, B 
                           => n3229, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128196792_128196960_128197184);
   U1590 : XOR2X1 port map( A => n411, B => n3231, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_127627392_128196680_128196848);
   U1591 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b12
                           , B => n3151, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831680_127845936_127847840);
   U1592 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b8,
                           B => n3145, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673568_127675472_127730688);
   U1593 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635920_127637824_127713520, B 
                           => n3217, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223888_128224112_128224056);
   U1594 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715536_127848576, B 
                           => n3223, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128224728_128224896_128225064);
   U1595 : OR3XL port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_3_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_4_port, C 
                           => n3813, Y => n3811);
   U1596 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_128223384_128223552);
   U1597 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_127826128_127826296);
   U1598 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263336_128263560_128263728, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263896_128264064_128264176, Y 
                           => n3304);
   U1599 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198864_128199032_128199200, B 
                           => n3282, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263896_128264064_128264176);
   U1600 : XOR2X1 port map( A => n399, B => n3281, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128263336_128263560_128263728);
   U1601 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127627504_127629408, B 
                           => n3244, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198864_128199032_128199200);
   U1602 : XOR2X1 port map( A => n400, B => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_17_port, Y 
                           => n2355);
   U1603 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128315744_128315968_128316136, B 
                           => n3324, Y => 
                           output_p1_times_a1_mul_componentxUMxsecond_vector_17_port);
   U1604 : INVX1 port map( A => n3323, Y => n400);
   U1605 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128237752_128237976_128238144, B 
                           => n3319, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer5_128315744_128315968_128316136);
   U1606 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128223384_128223552);
   U1607 : INVX1 port map( A => n4553, Y => n503);
   U1608 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_4_port, 
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_4_port, 
                           B1 => n4548, Y => n4553);
   U1609 : XOR2X1 port map( A => n3812, B => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_4_port, Y 
                           => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_4_port);
   U1610 : OR2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_3_port, B 
                           => n3813, Y => n3812);
   U1611 : INVX1 port map( A => n4551, Y => n488);
   U1612 : AOI22XL port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_6_port, 
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_6_port, 
                           B1 => n4548, Y => n4551);
   U1613 : XOR2X1 port map( A => n3810, B => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_6_port, Y 
                           => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_6_port);
   U1614 : OR2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_5_port, B 
                           => n3811, Y => n3810);
   U1615 : INVX1 port map( A => n3164, Y => n403);
   U1616 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b11, A1 
                           => output_p1_times_a1_mul_componentxUMxa3_and_b12, 
                           B0 => n3163, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b10, Y =>
                           n3164);
   U1617 : INVX1 port map( A => n3152, Y => n443);
   U1618 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b13, A1 
                           => output_p1_times_a1_mul_componentxUMxa0_and_b14, 
                           B0 => n3151, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b12, Y =>
                           n3152);
   U1619 : INVX1 port map( A => n3220, Y => n427);
   U1620 : AOI22X1 port map( A0 => n455, A1 => n428, B0 => n3219, B1 => n485, Y
                           => n3220);
   U1621 : INVX1 port map( A => n3270, Y => n419);
   U1622 : AOI22X1 port map( A0 => n427, A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
                           B0 => n3269, B1 => n420, Y => n3270);
   U1623 : AOI22X1 port map( A0 => output_previous_1_14_port, A1 => n133, B0 =>
                           output_p1_times_a1_mul_componentxinput_A_inverted_14_port, 
                           B1 => n165, Y => n4541);
   U1624 : XOR2X1 port map( A => n3787, B => output_previous_1_14_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_14_port);
   U1625 : OR2X2 port map( A => output_previous_1_13_port, B => n3786, Y => 
                           n3787);
   U1626 : INVX1 port map( A => n3162, Y => n444);
   U1627 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b14, A1 
                           => output_p1_times_a1_mul_componentxUMxa0_and_b15, 
                           B0 => n3161, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b13, Y =>
                           n3162);
   U1628 : INVX1 port map( A => n3224, Y => n475);
   U1629 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
                           B0 => n3223, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715536_127848576, Y 
                           => n3224);
   U1630 : INVX1 port map( A => n3226, Y => n424);
   U1631 : AOI22X1 port map( A0 => n446, A1 => n426, B0 => n3225, B1 => n474, Y
                           => n3226);
   U1632 : INVX1 port map( A => n3154, Y => n411);
   U1633 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b10, A1 
                           => output_p1_times_a1_mul_componentxUMxa3_and_b11, 
                           B0 => n3153, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b9, Y => 
                           n3154);
   U1634 : INVX1 port map( A => n3222, Y => n420);
   U1635 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
                           A1 => n504, B0 => n3221, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673568_127675472_127730688, Y 
                           => n3222);
   U1636 : INVX1 port map( A => n3230, Y => n413);
   U1637 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
                           B0 => n3229, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636144_127638048_127713744, Y 
                           => n3230);
   U1638 : AOI22X1 port map( A0 => output_previous_1_15_port, A1 => n133, B0 =>
                           output_p1_times_a1_mul_componentxinput_A_inverted_15_port, 
                           B1 => n165, Y => n4540);
   U1639 : XNOR2X1 port map( A => n3785, B => output_previous_1_15_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_15_port);
   U1640 : AOI22X1 port map( A0 => output_previous_1_16_port, A1 => n133, B0 =>
                           output_p1_times_a1_mul_componentxinput_A_inverted_16_port, 
                           B1 => n165, Y => n4539);
   U1641 : XNOR2X1 port map( A => n3784, B => output_previous_1_16_port, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_16_port);
   U1642 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b9, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b10, B0 
                           => n3175, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b8, Y => 
                           n3176);
   U1643 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b12, A1 
                           => output_p1_times_a1_mul_componentxUMxa3_and_b13, 
                           B0 => n3173, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b11, Y =>
                           n3174);
   U1644 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b8,
                           B => n3175, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732928_127722608_127724512);
   U1645 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b10
                           , B => output_p1_times_a1_mul_componentxUMxa7_and_b9
                           , Y => n3175);
   U1646 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b13
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b12, Y =>
                           n3173);
   U1647 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b16
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b15, Y =>
                           n3171);
   U1648 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b9,
                           B => output_p1_times_a1_mul_componentxUMxa7_and_b8, 
                           Y => n3165);
   U1649 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b11
                           , B => n3173, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673904_127675808_127731024);
   U1650 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198024_128197968);
   U1651 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b14
                           , B => n3171, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831904_127846160_127848064);
   U1652 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b7,
                           B => n3165, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732816_127722496_127724400);
   U1653 : OR3XL port map( A => n517, B => n516, C => n518, Y => n4003);
   U1654 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636368_127638272_127713968, B 
                           => n3241, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198472_128198640_128198808);
   U1655 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_128198024_128197968);
   U1656 : INVX1 port map( A => n4554, Y => n509);
   U1657 : AOI22XL port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_3_port, 
                           A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_3_port, 
                           B1 => n4548, Y => n4554);
   U1658 : XOR2X1 port map( A => n3813, B => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_3_port, Y 
                           => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_3_port);
   U1659 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_128198976_128199144, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198304_128198528_128198696, Y 
                           => n3282);
   U1660 : AND2X2 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer2_128198976_128199144);
   U1661 : XOR2X1 port map( A => n445, B => n3243, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198304_128198528_128198696);
   U1662 : INVX1 port map( A => n3176, Y => n445);
   U1663 : XOR2X1 port map( A => n3172, B => n3174, Y => n3243);
   U1664 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b15, A1 
                           => output_p1_times_a1_mul_componentxUMxa0_and_b16, 
                           B0 => n3171, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b14, Y =>
                           n3172);
   U1665 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128198976_128199144);
   U1666 : INVX1 port map( A => n3166, Y => n454);
   U1667 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b8, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b9, B0 =>
                           n3165, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b7, Y => 
                           n3166);
   U1668 : INVX1 port map( A => n3242, Y => n399);
   U1669 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
                           A1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
                           B0 => n3241, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636368_127638272_127713968, Y 
                           => n3242);
   U1670 : INVX1 port map( A => n3278, Y => n404);
   U1671 : AOI22X1 port map( A0 => n465, A1 => n410, B0 => n3277, B1 => n406, Y
                           => n3278);
   U1672 : XOR2X1 port map( A => n3783, B => n165, Y => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_17_port);
   U1673 : NAND2BX1 port map( AN => output_previous_1_16_port, B => n3784, Y =>
                           n3783);
   U1674 : XNOR2X1 port map( A => n516, B => n4004, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_2_port);
   U1675 : NOR2X1 port map( A => n518, B => n517, Y => n4004);
   U1676 : INVX1 port map( A => n3032, Y => n1068);
   U1677 : AOI22X1 port map( A0 => n1069, A1 => n1070, B0 => n3031, B1 => n1092
                           , Y => n3032);
   U1678 : INVX1 port map( A => n3500, Y => n591);
   U1679 : AOI22X1 port map( A0 => n592, A1 => n593, B0 => n3499, B1 => n615, Y
                           => n3500);
   U1680 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831456_127845712_127847616, B 
                           => n2747, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223440_128223608_128223776);
   U1681 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831456_127845712_127847616, B 
                           => n2981, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223440_128223608_128223776);
   U1682 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831456_127845712_127847616, B 
                           => n3449, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223440_128223608_128223776);
   U1683 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831456_127845712_127847616, B 
                           => n2513, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223440_128223608_128223776);
   U1684 : XOR2X1 port map( A => n968, B => n988, Y => n2747);
   U1685 : XOR2X1 port map( A => n1127, B => n1147, Y => n2981);
   U1686 : XOR2X1 port map( A => n650, B => n670, Y => n3449);
   U1687 : XOR2X1 port map( A => n809, B => n829, Y => n2513);
   U1688 : XOR2X1 port map( A => n911, B => n910, Y => n2797);
   U1689 : XOR2X1 port map( A => n1070, B => n1069, Y => n3031);
   U1690 : XOR2X1 port map( A => n593, B => n592, Y => n3499);
   U1691 : XOR2X1 port map( A => n752, B => n751, Y => n2563);
   U1692 : BUFX3 port map( A => n4451, Y => n190);
   U1693 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_17, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_17_port, 
                           B1 => n4442, Y => n4451);
   U1694 : XOR2X1 port map( A => n3719, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_17, 
                           Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_17_port);
   U1695 : XOR2X1 port map( A => n2312, B => n2313, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_17);
   U1696 : BUFX3 port map( A => n4504, Y => n211);
   U1697 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_17, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_17_port, 
                           B1 => n4495, Y => n4504);
   U1698 : XOR2X1 port map( A => n3767, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_17, 
                           Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_17_port);
   U1699 : XOR2X1 port map( A => n2333, B => n2334, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_17);
   U1700 : BUFX3 port map( A => n4610, Y => n253);
   U1701 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_17,
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_17_port, 
                           B1 => n4601, Y => n4610);
   U1702 : XOR2X1 port map( A => n3863, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_17,
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_17_port);
   U1703 : XOR2X1 port map( A => n2375, B => n2376, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_17)
                           ;
   U1704 : BUFX3 port map( A => input_times_b0_mul_componentxn100, Y => n281);
   U1705 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_17, A1 
                           => n121, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_17_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn100);
   U1706 : XOR2X1 port map( A => n3671, B => 
                           input_times_b0_mul_componentxunsigned_output_17, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_17_port);
   U1707 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxAdder_finalxn474, B 
                           => input_times_b0_mul_componentxUMxAdder_finalxn475,
                           Y => input_times_b0_mul_componentxunsigned_output_17
                           );
   U1708 : INVX1 port map( A => n2748, Y => n910);
   U1709 : AOI22X1 port map( A0 => n988, A1 => n968, B0 => n2747, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831456_127845712_127847616, Y 
                           => n2748);
   U1710 : INVX1 port map( A => n2982, Y => n1069);
   U1711 : AOI22X1 port map( A0 => n1147, A1 => n1127, B0 => n2981, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831456_127845712_127847616, Y 
                           => n2982);
   U1712 : INVX1 port map( A => n3450, Y => n592);
   U1713 : AOI22X1 port map( A0 => n670, A1 => n650, B0 => n3449, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831456_127845712_127847616, Y 
                           => n3450);
   U1714 : INVX1 port map( A => n2514, Y => n751);
   U1715 : AOI22X1 port map( A0 => n829, A1 => n809, B0 => n2513, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831456_127845712_127847616, Y 
                           => n2514);
   U1716 : INVX1 port map( A => n2798, Y => n909);
   U1717 : AOI22X1 port map( A0 => n910, A1 => n911, B0 => n2797, B1 => n933, Y
                           => n2798);
   U1718 : INVX1 port map( A => n2564, Y => n750);
   U1719 : AOI22X1 port map( A0 => n751, A1 => n752, B0 => n2563, B1 => n774, Y
                           => n2564);
   U1720 : XOR2X1 port map( A => n517, B => n518, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_1_port);
   U1721 : INVX1 port map( A => n4510, Y => n1076);
   U1722 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_11, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_11_port, 
                           B1 => n4495, Y => n4510);
   U1723 : XOR2X1 port map( A => n3772, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_11, 
                           Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_11_port);
   U1724 : INVX1 port map( A => n4616, Y => n599);
   U1725 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_11,
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_11_port, 
                           B1 => n4601, Y => n4616);
   U1726 : XOR2X1 port map( A => n3868, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_11,
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_11_port);
   U1727 : INVX1 port map( A => n2722, Y => n979);
   U1728 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
                           A1 => n985, B0 => n2721, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672560_127674464, Y 
                           => n2722);
   U1729 : INVX1 port map( A => n2956, Y => n1138);
   U1730 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
                           A1 => n1144, B0 => n2955, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672560_127674464, Y 
                           => n2956);
   U1731 : INVX1 port map( A => n3424, Y => n661);
   U1732 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
                           A1 => n667, B0 => n3423, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672560_127674464, Y 
                           => n3424);
   U1733 : INVX1 port map( A => n2488, Y => n820);
   U1734 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830560_127844816_127846720, 
                           A1 => n826, B0 => n2487, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672560_127674464, Y 
                           => n2488);
   U1735 : INVX1 port map( A => n2974, Y => n1087);
   U1736 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
                           B0 => n2973, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732256_127721936_127723840, Y 
                           => n2974);
   U1737 : INVX1 port map( A => n3442, Y => n610);
   U1738 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
                           B0 => n3441, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732256_127721936_127723840, Y 
                           => n3442);
   U1739 : INVX1 port map( A => n2756, Y => n952);
   U1740 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
                           B0 => n2755, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715536_127848576, Y 
                           => n2756);
   U1741 : INVX1 port map( A => n2978, Y => n1074);
   U1742 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127635696_127637600, 
                           B0 => n2977, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673344_127675248_127730464, Y 
                           => n2978);
   U1743 : INVX1 port map( A => n3446, Y => n597);
   U1744 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127635696_127637600, 
                           B0 => n3445, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673344_127675248_127730464, Y 
                           => n3446);
   U1745 : INVX1 port map( A => n2522, Y => n793);
   U1746 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
                           B0 => n2521, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715536_127848576, Y 
                           => n2522);
   U1747 : AOI22X1 port map( A0 => n984, A1 => n961, B0 => n2771, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831904_127846160_127848064, Y 
                           => n2772);
   U1748 : AOI22X1 port map( A0 => n1143, A1 => n1120, B0 => n3005, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831904_127846160_127848064, Y 
                           => n3006);
   U1749 : AOI22X1 port map( A0 => n666, A1 => n643, B0 => n3473, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831904_127846160_127848064, Y 
                           => n3474);
   U1750 : AOI22X1 port map( A0 => n825, A1 => n802, B0 => n2537, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831904_127846160_127848064, Y 
                           => n2538);
   U1751 : INVX1 port map( A => n2738, Y => n934);
   U1752 : AOI22X1 port map( A0 => n963, A1 => n935, B0 => n2737, B1 => n982, Y
                           => n2738);
   U1753 : INVX1 port map( A => n2972, Y => n1093);
   U1754 : AOI22X1 port map( A0 => n1122, A1 => n1094, B0 => n2971, B1 => n1141
                           , Y => n2972);
   U1755 : INVX1 port map( A => n3440, Y => n616);
   U1756 : AOI22X1 port map( A0 => n645, A1 => n617, B0 => n3439, B1 => n664, Y
                           => n3440);
   U1757 : INVX1 port map( A => n2504, Y => n775);
   U1758 : AOI22X1 port map( A0 => n804, A1 => n776, B0 => n2503, B1 => n823, Y
                           => n2504);
   U1759 : INVX1 port map( A => n3022, Y => n1106);
   U1760 : AOI22X1 port map( A0 => n1113, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
                           B0 => n3021, B1 => n1107, Y => n3022);
   U1761 : INVX1 port map( A => n3490, Y => n629);
   U1762 : AOI22X1 port map( A0 => n636, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
                           B0 => n3489, B1 => n630, Y => n3490);
   U1763 : INVX1 port map( A => n2742, Y => n924);
   U1764 : AOI22X1 port map( A0 => n953, A1 => n927, B0 => n2741, B1 => n976, Y
                           => n2742);
   U1765 : INVX1 port map( A => n2508, Y => n765);
   U1766 : AOI22X1 port map( A0 => n794, A1 => n768, B0 => n2507, B1 => n817, Y
                           => n2508);
   U1767 : XOR2X1 port map( A => n990, B => n2725, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127731808_127826912_127827136);
   U1768 : XOR2X1 port map( A => n1149, B => n2959, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127731808_127826912_127827136);
   U1769 : XOR2X1 port map( A => n672, B => n3427, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127731808_127826912_127827136);
   U1770 : XOR2X1 port map( A => n831, B => n2491, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127731808_127826912_127827136);
   U1771 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673568_127675472_127730688, B 
                           => n2753, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224280_128224448_128224560);
   U1772 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673568_127675472_127730688, B 
                           => n2987, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224280_128224448_128224560);
   U1773 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673568_127675472_127730688, B 
                           => n3455, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224280_128224448_128224560);
   U1774 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673568_127675472_127730688, B 
                           => n2519, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224280_128224448_128224560);
   U1775 : XOR2X1 port map( A => n991, B => n2765, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197016_128197240_128197352);
   U1776 : XOR2X1 port map( A => n1150, B => n2999, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197016_128197240_128197352);
   U1777 : XOR2X1 port map( A => n673, B => n3467, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197016_128197240_128197352);
   U1778 : XOR2X1 port map( A => n832, B => n2531, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197016_128197240_128197352);
   U1779 : XOR2X1 port map( A => n978, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127672560_127674464, Y 
                           => n2723);
   U1780 : XOR2X1 port map( A => n1137, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127672560_127674464, Y 
                           => n2957);
   U1781 : XOR2X1 port map( A => n660, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127672560_127674464, Y 
                           => n3425);
   U1782 : XOR2X1 port map( A => n819, B => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127672560_127674464, Y 
                           => n2489);
   U1783 : XOR2X1 port map( A => n985, B => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830560_127844816_127846720, Y 
                           => n2721);
   U1784 : XOR2X1 port map( A => n1144, B => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830560_127844816_127846720, Y 
                           => n2955);
   U1785 : XOR2X1 port map( A => n667, B => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830560_127844816_127846720, Y 
                           => n3423);
   U1786 : XOR2X1 port map( A => n826, B => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830560_127844816_127846720, Y 
                           => n2487);
   U1787 : XOR2X1 port map( A => n970, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127827304_127827416, Y 
                           => n2783);
   U1788 : XOR2X1 port map( A => n989, B => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831120_127845376_127847280, Y 
                           => n2735);
   U1789 : XOR2X1 port map( A => n1129, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127827304_127827416, Y 
                           => n3017);
   U1790 : XOR2X1 port map( A => n1148, B => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831120_127845376_127847280, Y 
                           => n2969);
   U1791 : XOR2X1 port map( A => n652, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127827304_127827416, Y 
                           => n3485);
   U1792 : XOR2X1 port map( A => n671, B => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831120_127845376_127847280, Y 
                           => n3437);
   U1793 : XOR2X1 port map( A => n811, B => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127827304_127827416, Y 
                           => n2549);
   U1794 : XOR2X1 port map( A => n830, B => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831120_127845376_127847280, Y 
                           => n2501);
   U1795 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831008_127845264_127847168, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673008_127674912_127730128, Y 
                           => n2731);
   U1796 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831008_127845264_127847168, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673008_127674912_127730128, Y 
                           => n2965);
   U1797 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831008_127845264_127847168, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673008_127674912_127730128, Y 
                           => n3433);
   U1798 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831008_127845264_127847168, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673008_127674912_127730128, Y 
                           => n2497);
   U1799 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831232_127845488_127847392, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673232_127675136_127730352, Y 
                           => n2739);
   U1800 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831232_127845488_127847392, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673232_127675136_127730352, Y 
                           => n2973);
   U1801 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831232_127845488_127847392, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673232_127675136_127730352, Y 
                           => n3441);
   U1802 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831232_127845488_127847392, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673232_127675136_127730352, Y 
                           => n2505);
   U1803 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673456_127675360_127730576, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732480_127722160_127724064, Y 
                           => n2749);
   U1804 : XOR2X1 port map( A => n981, B => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831568_127845824_127847728, Y 
                           => n2753);
   U1805 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732592_127722272_127724176, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636032_127637936_127713632, Y 
                           => n2755);
   U1806 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673456_127675360_127730576, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732480_127722160_127724064, Y 
                           => n2983);
   U1807 : XOR2X1 port map( A => n1140, B => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831568_127845824_127847728, Y 
                           => n2987);
   U1808 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732592_127722272_127724176, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636032_127637936_127713632, Y 
                           => n2989);
   U1809 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673456_127675360_127730576, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732480_127722160_127724064, Y 
                           => n3451);
   U1810 : XOR2X1 port map( A => n663, B => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831568_127845824_127847728, Y 
                           => n3455);
   U1811 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732592_127722272_127724176, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636032_127637936_127713632, Y 
                           => n3457);
   U1812 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673456_127675360_127730576, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732480_127722160_127724064, Y 
                           => n2515);
   U1813 : XOR2X1 port map( A => n822, B => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831568_127845824_127847728, Y 
                           => n2519);
   U1814 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732592_127722272_127724176, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636032_127637936_127713632, Y 
                           => n2521);
   U1815 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127635696_127637600, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831344_127845600_127847504, Y 
                           => n2743);
   U1816 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127635696_127637600, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831344_127845600_127847504, Y 
                           => n2977);
   U1817 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127635696_127637600, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831344_127845600_127847504, Y 
                           => n3445);
   U1818 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127635696_127637600, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831344_127845600_127847504, Y 
                           => n2509);
   U1819 : XOR2X1 port map( A => n975, B => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127715536_127848576, Y 
                           => n2759);
   U1820 : XOR2X1 port map( A => n1134, B => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127715536_127848576, Y 
                           => n2993);
   U1821 : XOR2X1 port map( A => n657, B => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127715536_127848576, Y 
                           => n3461);
   U1822 : XOR2X1 port map( A => n816, B => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127715536_127848576, Y 
                           => n2525);
   U1823 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673680_127675584_127730800, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732704_127722384_127724288, Y 
                           => n2761);
   U1824 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673680_127675584_127730800, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732704_127722384_127724288, Y 
                           => n2527);
   U1825 : XOR2X1 port map( A => n964, B => n983, Y => n2727);
   U1826 : XOR2X1 port map( A => n956, B => n977, Y => n2729);
   U1827 : XOR2X1 port map( A => n1123, B => n1142, Y => n2961);
   U1828 : XOR2X1 port map( A => n1115, B => n1136, Y => n2963);
   U1829 : XOR2X1 port map( A => n646, B => n665, Y => n3429);
   U1830 : XOR2X1 port map( A => n638, B => n659, Y => n3431);
   U1831 : XOR2X1 port map( A => n805, B => n824, Y => n2493);
   U1832 : XOR2X1 port map( A => n797, B => n818, Y => n2495);
   U1833 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672672_127674576_127729792, B 
                           => n979, Y => n2779);
   U1834 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672672_127674576_127729792, B 
                           => n1138, Y => n3013);
   U1835 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672672_127674576_127729792, B 
                           => n661, Y => n3481);
   U1836 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672672_127674576_127729792, B 
                           => n820, Y => n2545);
   U1837 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635696_127637600, B 
                           => n945, Y => n2789);
   U1838 : XOR2X1 port map( A => n935, B => n963, Y => n2737);
   U1839 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732144_127721824_127723728, B 
                           => n954, Y => n2787);
   U1840 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635696_127637600, B 
                           => n1104, Y => n3023);
   U1841 : XOR2X1 port map( A => n1094, B => n1122, Y => n2971);
   U1842 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732144_127721824_127723728, B 
                           => n1113, Y => n3021);
   U1843 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635696_127637600, B 
                           => n627, Y => n3491);
   U1844 : XOR2X1 port map( A => n617, B => n645, Y => n3439);
   U1845 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732144_127721824_127723728, B 
                           => n636, Y => n3489);
   U1846 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635696_127637600, B 
                           => n786, Y => n2555);
   U1847 : XOR2X1 port map( A => n776, B => n804, Y => n2503);
   U1848 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732144_127721824_127723728, B 
                           => n795, Y => n2553);
   U1849 : XOR2X1 port map( A => n927, B => n953, Y => n2741);
   U1850 : XOR2X1 port map( A => n1086, B => n1112, Y => n2975);
   U1851 : XOR2X1 port map( A => n609, B => n635, Y => n3443);
   U1852 : XOR2X1 port map( A => n768, B => n794, Y => n2507);
   U1853 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715648_127848688_127850592, B 
                           => n903, Y => n2801);
   U1854 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715648_127848688_127850592, B 
                           => n1062, Y => n3035);
   U1855 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715648_127848688_127850592, B 
                           => n585, Y => n3503);
   U1856 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715648_127848688_127850592, B 
                           => n744, Y => n2567);
   U1857 : XOR2X1 port map( A => n943, B => n967, Y => n2765);
   U1858 : XOR2X1 port map( A => n1102, B => n1126, Y => n2999);
   U1859 : XOR2X1 port map( A => n625, B => n649, Y => n3467);
   U1860 : XOR2X1 port map( A => n784, B => n808, Y => n2531);
   U1861 : XOR2X1 port map( A => n961, B => n984, Y => n2771);
   U1862 : XOR2X1 port map( A => n1120, B => n1143, Y => n3005);
   U1863 : XOR2X1 port map( A => n643, B => n666, Y => n3473);
   U1864 : XOR2X1 port map( A => n802, B => n825, Y => n2537);
   U1865 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127827304_127827416);
   U1866 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127827304_127827416);
   U1867 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127827304_127827416);
   U1868 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127827304_127827416);
   U1869 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127827752_127827920);
   U1870 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127827752_127827920);
   U1871 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127827752_127827920);
   U1872 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127827752_127827920);
   U1873 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827752_127827920);
   U1874 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827752_127827920);
   U1875 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732032_127721712_127723616, B 
                           => n2731, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221424_128221536_128221704);
   U1876 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732032_127721712_127723616, B 
                           => n2965, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221424_128221536_128221704);
   U1877 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732032_127721712_127723616, B 
                           => n3433, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221424_128221536_128221704);
   U1878 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732032_127721712_127723616, B 
                           => n2497, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221424_128221536_128221704);
   U1879 : XOR2X1 port map( A => n944, B => n2745, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127715424_128223048_128223272);
   U1880 : XOR2X1 port map( A => n1103, B => n2979, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127715424_128223048_128223272);
   U1881 : XOR2X1 port map( A => n626, B => n3447, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127715424_128223048_128223272);
   U1882 : XOR2X1 port map( A => n785, B => n2511, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127715424_128223048_128223272);
   U1883 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636144_127638048_127713744, B 
                           => n2761, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128196792_128196960_128197184);
   U1884 : XOR2X1 port map( A => n887, B => n2763, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127627392_128196680_128196848);
   U1885 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636144_127638048_127713744, B 
                           => n2995, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128196792_128196960_128197184);
   U1886 : XOR2X1 port map( A => n1046, B => n2997, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127627392_128196680_128196848);
   U1887 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636144_127638048_127713744, B 
                           => n3463, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128196792_128196960_128197184);
   U1888 : XOR2X1 port map( A => n569, B => n3465, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127627392_128196680_128196848);
   U1889 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636144_127638048_127713744, B 
                           => n2527, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128196792_128196960_128197184);
   U1890 : XOR2X1 port map( A => n728, B => n2529, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127627392_128196680_128196848);
   U1891 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827304_127827416);
   U1892 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827304_127827416);
   U1893 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827304_127827416);
   U1894 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672784_127674688_127729904, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830784_127845040_127846944, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827304_127827416);
   U1895 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830896_127845152_127847056, B 
                           => n2727, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827248_127827472_127827640);
   U1896 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830896_127845152_127847056, B 
                           => n2961, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827248_127827472_127827640);
   U1897 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830896_127845152_127847056, B 
                           => n3429, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827248_127827472_127827640);
   U1898 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830896_127845152_127847056, B 
                           => n2493, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827248_127827472_127827640);
   U1899 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127731920_127721600, B 
                           => n2729, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827584_127827808_128221256);
   U1900 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127731920_127721600, B 
                           => n2963, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827584_127827808_128221256);
   U1901 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127731920_127721600, B 
                           => n3431, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827584_127827808_128221256);
   U1902 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127731920_127721600, B 
                           => n2495, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827584_127827808_128221256);
   U1903 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635920_127637824_127713520, B 
                           => n2749, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223888_128224112_128224056);
   U1904 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831680_127845936_127847840, B 
                           => n2759, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224952_128225120_128225232);
   U1905 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635920_127637824_127713520, B 
                           => n2983, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223888_128224112_128224056);
   U1906 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831680_127845936_127847840, B 
                           => n2993, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224952_128225120_128225232);
   U1907 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635920_127637824_127713520, B 
                           => n3451, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223888_128224112_128224056);
   U1908 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831680_127845936_127847840, B 
                           => n3461, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224952_128225120_128225232);
   U1909 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635920_127637824_127713520, B 
                           => n2515, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223888_128224112_128224056);
   U1910 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831680_127845936_127847840, B 
                           => n2525, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224952_128225120_128225232);
   U1911 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715536_127848576, B 
                           => n2755, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224728_128224896_128225064);
   U1912 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715536_127848576, B 
                           => n2989, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224728_128224896_128225064);
   U1913 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715536_127848576, B 
                           => n3457, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224728_128224896_128225064);
   U1914 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715536_127848576, B 
                           => n2521, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224728_128224896_128225064);
   U1915 : XOR2X1 port map( A => n982, B => n2737, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221872_128222096_128222264);
   U1916 : XOR2X1 port map( A => n969, B => n2733, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127635584_128221368_128221592);
   U1917 : XOR2X1 port map( A => n1141, B => n2971, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221872_128222096_128222264);
   U1918 : XOR2X1 port map( A => n1128, B => n2967, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127635584_128221368_128221592);
   U1919 : XOR2X1 port map( A => n664, B => n3439, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221872_128222096_128222264);
   U1920 : XOR2X1 port map( A => n651, B => n3435, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127635584_128221368_128221592);
   U1921 : XOR2X1 port map( A => n823, B => n2503, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221872_128222096_128222264);
   U1922 : XOR2X1 port map( A => n810, B => n2499, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127635584_128221368_128221592);
   U1923 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673344_127675248_127730464, B 
                           => n2743, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222936_128223104_128223216);
   U1924 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673344_127675248_127730464, B 
                           => n2977, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222936_128223104_128223216);
   U1925 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673344_127675248_127730464, B 
                           => n3445, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222936_128223104_128223216);
   U1926 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673344_127675248_127730464, B 
                           => n2509, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222936_128223104_128223216);
   U1927 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_128223384_128223552);
   U1928 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_128223384_128223552);
   U1929 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_128223384_128223552);
   U1930 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer2_128223384_128223552);
   U1931 : INVX1 port map( A => n4455, Y => n899);
   U1932 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_13, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_13_port, 
                           B1 => n4442, Y => n4455);
   U1933 : XOR2X1 port map( A => n3722, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_13, 
                           Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_13_port);
   U1934 : INVX1 port map( A => n4508, Y => n1058);
   U1935 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_13, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_13_port, 
                           B1 => n4495, Y => n4508);
   U1936 : XOR2X1 port map( A => n3770, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_13, 
                           Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_13_port);
   U1937 : INVX1 port map( A => n4614, Y => n581);
   U1938 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_13,
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_13_port, 
                           B1 => n4601, Y => n4614);
   U1939 : XOR2X1 port map( A => n3866, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_13,
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_13_port);
   U1940 : INVX1 port map( A => input_times_b0_mul_componentxn104, Y => n740);
   U1941 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_13, A1 
                           => n121, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_13_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn104);
   U1942 : XOR2X1 port map( A => n3674, B => 
                           input_times_b0_mul_componentxunsigned_output_13, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_13_port);
   U1943 : INVX1 port map( A => n4453, Y => n884);
   U1944 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_15, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_15_port, 
                           B1 => n4442, Y => n4453);
   U1945 : XNOR2X1 port map( A => n3721, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_15, 
                           Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_15_port);
   U1946 : INVX1 port map( A => input_times_b0_mul_componentxn102, Y => n725);
   U1947 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_15, A1 
                           => n121, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_15_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn102);
   U1948 : XNOR2X1 port map( A => n3673, B => 
                           input_times_b0_mul_componentxunsigned_output_15, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_15_port);
   U1949 : INVX1 port map( A => n4454, Y => n893);
   U1950 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_14, 
                           A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_14_port, 
                           B1 => n4442, Y => n4454);
   U1951 : XOR2X1 port map( A => n3723, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_14, 
                           Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_14_port);
   U1952 : OR2X2 port map( A => 
                           input_p1_times_b1_mul_componentxunsigned_output_13, 
                           B => n3722, Y => n3723);
   U1953 : INVX1 port map( A => n4507, Y => n1052);
   U1954 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_14, 
                           A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_14_port, 
                           B1 => n4495, Y => n4507);
   U1955 : XOR2X1 port map( A => n3771, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_14, 
                           Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_14_port);
   U1956 : OR2X2 port map( A => 
                           input_p2_times_b2_mul_componentxunsigned_output_13, 
                           B => n3770, Y => n3771);
   U1957 : INVX1 port map( A => n4613, Y => n575);
   U1958 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_14,
                           A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_14_port, 
                           B1 => n4601, Y => n4613);
   U1959 : XOR2X1 port map( A => n3867, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_14,
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_14_port);
   U1960 : OR2X2 port map( A => 
                           output_p2_times_a2_mul_componentxunsigned_output_13,
                           B => n3866, Y => n3867);
   U1961 : INVX1 port map( A => input_times_b0_mul_componentxn103, Y => n734);
   U1962 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_14, A1 
                           => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_14_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn103);
   U1963 : XOR2X1 port map( A => n3675, B => 
                           input_times_b0_mul_componentxunsigned_output_14, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_14_port);
   U1964 : OR2X2 port map( A => input_times_b0_mul_componentxunsigned_output_13
                           , B => n3674, Y => n3675);
   U1965 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263336_128263560_128263728, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263896_128264064_128264176, Y 
                           => n2836);
   U1966 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198864_128199032_128199200, B 
                           => n2814, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263896_128264064_128264176);
   U1967 : XOR2X1 port map( A => n874, B => n2813, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128263336_128263560_128263728);
   U1968 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127627504_127629408, B 
                           => n2776, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198864_128199032_128199200);
   U1969 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263336_128263560_128263728, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263896_128264064_128264176, Y 
                           => n3070);
   U1970 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198864_128199032_128199200, B 
                           => n3048, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263896_128264064_128264176);
   U1971 : XOR2X1 port map( A => n1033, B => n3047, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128263336_128263560_128263728);
   U1972 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127627504_127629408, B 
                           => n3010, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198864_128199032_128199200);
   U1973 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263336_128263560_128263728, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263896_128264064_128264176, Y 
                           => n3538);
   U1974 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198864_128199032_128199200, B 
                           => n3516, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263896_128264064_128264176);
   U1975 : XOR2X1 port map( A => n556, B => n3515, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128263336_128263560_128263728);
   U1976 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127627504_127629408, B 
                           => n3478, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198864_128199032_128199200);
   U1977 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263336_128263560_128263728, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263896_128264064_128264176, Y 
                           => n2602);
   U1978 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198864_128199032_128199200, B 
                           => n2580, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263896_128264064_128264176);
   U1979 : XOR2X1 port map( A => n715, B => n2579, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128263336_128263560_128263728);
   U1980 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127627504_127629408, B 
                           => n2542, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198864_128199032_128199200);
   U1981 : XOR2X1 port map( A => n2770, B => n2772, Y => n2813);
   U1982 : AOI22X1 port map( A0 => n879, A1 => n920, B0 => n2769, B1 => n931, Y
                           => n2770);
   U1983 : XOR2X1 port map( A => n3004, B => n3006, Y => n3047);
   U1984 : AOI22X1 port map( A0 => n1038, A1 => n1079, B0 => n3003, B1 => n1090
                           , Y => n3004);
   U1985 : XOR2X1 port map( A => n3472, B => n3474, Y => n3515);
   U1986 : AOI22X1 port map( A0 => n561, A1 => n602, B0 => n3471, B1 => n613, Y
                           => n3472);
   U1987 : XOR2X1 port map( A => n2536, B => n2538, Y => n2579);
   U1988 : AOI22X1 port map( A0 => n720, A1 => n761, B0 => n2535, B1 => n772, Y
                           => n2536);
   U1989 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128238312_128238424_128238592, B 
                           => n881, Y => n2856);
   U1990 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128264344_128264512, B 
                           => n2836, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer4_128238312_128238424_128238592);
   U1991 : INVX1 port map( A => n2850, Y => n881);
   U1992 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128199816_128200040_128199984, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128199368_128199480_128199648, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128264344_128264512);
   U1993 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128238312_128238424_128238592, B 
                           => n1040, Y => n3090);
   U1994 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128264344_128264512, B 
                           => n3070, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer4_128238312_128238424_128238592);
   U1995 : INVX1 port map( A => n3084, Y => n1040);
   U1996 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128199816_128200040_128199984, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128199368_128199480_128199648, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128264344_128264512);
   U1997 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128238312_128238424_128238592, B 
                           => n563, Y => n3558);
   U1998 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128264344_128264512, B 
                           => n3538, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer4_128238312_128238424_128238592);
   U1999 : INVX1 port map( A => n3552, Y => n563);
   U2000 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128199816_128200040_128199984, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128199368_128199480_128199648, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128264344_128264512);
   U2001 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer4_128238312_128238424_128238592, B 
                           => n722, Y => n2622);
   U2002 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer3_128264344_128264512, B 
                           => n2602, Y => 
                           input_times_b0_mul_componentxUMxsum_layer4_128238312_128238424_128238592);
   U2003 : INVX1 port map( A => n2616, Y => n722);
   U2004 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_128199816_128200040_128199984, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128199368_128199480_128199648, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer3_128264344_128264512);
   U2005 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223384_128223552);
   U2006 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223384_128223552);
   U2007 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223384_128223552);
   U2008 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635808_127637712_127713408, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732368_127722048_127723952, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223384_128223552);
   U2009 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732256_127721936_127723840, B 
                           => n2739, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222432_128222544_128222712);
   U2010 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673120_127675024_127730240, B 
                           => n2735, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128221760_128221928_128222040);
   U2011 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732256_127721936_127723840, B 
                           => n2973, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222432_128222544_128222712);
   U2012 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673120_127675024_127730240, B 
                           => n2969, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128221760_128221928_128222040);
   U2013 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732256_127721936_127723840, B 
                           => n3441, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222432_128222544_128222712);
   U2014 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673120_127675024_127730240, B 
                           => n3437, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128221760_128221928_128222040);
   U2015 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732256_127721936_127723840, B 
                           => n2505, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222432_128222544_128222712);
   U2016 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673120_127675024_127730240, B 
                           => n2501, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128221760_128221928_128222040);
   U2017 : INVX1 port map( A => n4456, Y => n908);
   U2018 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_12, 
                           A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_12_port, 
                           B1 => n4442, Y => n4456);
   U2019 : XOR2X1 port map( A => n3725, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_12, 
                           Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_12_port);
   U2020 : OR2X2 port map( A => n3724, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_11, 
                           Y => n3725);
   U2021 : INVX1 port map( A => n4509, Y => n1067);
   U2022 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_12, 
                           A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_12_port, 
                           B1 => n4495, Y => n4509);
   U2023 : XOR2X1 port map( A => n3773, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_12, 
                           Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_12_port);
   U2024 : OR2X2 port map( A => n3772, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_11, 
                           Y => n3773);
   U2025 : INVX1 port map( A => n4615, Y => n590);
   U2026 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_12,
                           A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_12_port, 
                           B1 => n4601, Y => n4615);
   U2027 : XOR2X1 port map( A => n3869, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_12,
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_12_port);
   U2028 : OR2X2 port map( A => n3868, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_11,
                           Y => n3869);
   U2029 : INVX1 port map( A => input_times_b0_mul_componentxn105, Y => n749);
   U2030 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_12, A1 
                           => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_12_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn105);
   U2031 : XOR2X1 port map( A => n3677, B => 
                           input_times_b0_mul_componentxunsigned_output_12, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_12_port);
   U2032 : OR2X2 port map( A => n3676, B => 
                           input_times_b0_mul_componentxunsigned_output_11, Y 
                           => n3677);
   U2033 : INVX1 port map( A => n4458, Y => n930);
   U2034 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_10, 
                           A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_10_port, 
                           B1 => n4442, Y => n4458);
   U2035 : XOR2X1 port map( A => n3726, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_10, 
                           Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_10_port);
   U2036 : NAND2X1 port map( A => n3711, B => n939, Y => n3726);
   U2037 : INVX1 port map( A => n4511, Y => n1089);
   U2038 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_10, 
                           A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_10_port, 
                           B1 => n4495, Y => n4511);
   U2039 : XOR2X1 port map( A => n3774, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_10, 
                           Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_10_port);
   U2040 : NAND2X1 port map( A => n3759, B => n1098, Y => n3774);
   U2041 : INVX1 port map( A => n4617, Y => n612);
   U2042 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_10,
                           A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_10_port, 
                           B1 => n4601, Y => n4617);
   U2043 : XOR2X1 port map( A => n3870, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_10,
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_10_port);
   U2044 : NAND2X1 port map( A => n3855, B => n621, Y => n3870);
   U2045 : INVX1 port map( A => input_times_b0_mul_componentxn107, Y => n771);
   U2046 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_10, A1 
                           => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_10_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn107);
   U2047 : XOR2X1 port map( A => n3678, B => 
                           input_times_b0_mul_componentxunsigned_output_10, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_10_port);
   U2048 : NAND2X1 port map( A => n3663, B => n780, Y => n3678);
   U2049 : INVX1 port map( A => n4452, Y => n876);
   U2050 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_16, 
                           A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_16_port, 
                           B1 => n4442, Y => n4452);
   U2051 : XNOR2X1 port map( A => n3720, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_16, 
                           Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_16_port);
   U2052 : INVX1 port map( A => input_times_b0_mul_componentxn101, Y => n717);
   U2053 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_16, A1 
                           => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_16_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn101);
   U2054 : XNOR2X1 port map( A => n3672, B => 
                           input_times_b0_mul_componentxunsigned_output_16, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_16_port);
   U2055 : INVX1 port map( A => n2730, Y => n954);
   U2056 : AOI22X1 port map( A0 => n977, A1 => n956, B0 => n2729, B1 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127731920_127721600, Y 
                           => n2730);
   U2057 : INVX1 port map( A => n2964, Y => n1113);
   U2058 : AOI22X1 port map( A0 => n1136, A1 => n1115, B0 => n2963, B1 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127731920_127721600, Y 
                           => n2964);
   U2059 : INVX1 port map( A => n3432, Y => n636);
   U2060 : AOI22X1 port map( A0 => n659, A1 => n638, B0 => n3431, B1 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127731920_127721600, Y 
                           => n3432);
   U2061 : INVX1 port map( A => n2496, Y => n795);
   U2062 : AOI22X1 port map( A0 => n818, A1 => n797, B0 => n2495, B1 => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127731920_127721600, Y 
                           => n2496);
   U2063 : INVX1 port map( A => n2784, Y => n959);
   U2064 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127827304_127827416, 
                           A1 => n970, B0 => n2783, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127827248_127827472_127827640, Y 
                           => n2784);
   U2065 : INVX1 port map( A => n3018, Y => n1118);
   U2066 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127827304_127827416, 
                           A1 => n1129, B0 => n3017, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827248_127827472_127827640, Y 
                           => n3018);
   U2067 : INVX1 port map( A => n3486, Y => n641);
   U2068 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127827304_127827416, 
                           A1 => n652, B0 => n3485, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827248_127827472_127827640, Y 
                           => n3486);
   U2069 : INVX1 port map( A => n2550, Y => n800);
   U2070 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127827304_127827416, 
                           A1 => n811, B0 => n2549, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_127827248_127827472_127827640, Y 
                           => n2550);
   U2071 : INVX1 port map( A => n2740, Y => n928);
   U2072 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
                           B0 => n2739, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732256_127721936_127723840, Y 
                           => n2740);
   U2073 : INVX1 port map( A => n2506, Y => n769);
   U2074 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673232_127675136_127730352, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831232_127845488_127847392, 
                           B0 => n2505, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732256_127721936_127723840, Y 
                           => n2506);
   U2075 : INVX1 port map( A => n2744, Y => n915);
   U2076 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127635696_127637600, 
                           B0 => n2743, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673344_127675248_127730464, Y 
                           => n2744);
   U2077 : INVX1 port map( A => n2510, Y => n756);
   U2078 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831344_127845600_127847504, 
                           A1 => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127635696_127637600, 
                           B0 => n2509, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673344_127675248_127730464, Y 
                           => n2510);
   U2079 : INVX1 port map( A => n2802, Y => n895);
   U2080 : AOI22X1 port map( A0 => n903, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
                           B0 => n2801, B1 => n896, Y => n2802);
   U2081 : INVX1 port map( A => n2760, Y => n918);
   U2082 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127715536_127848576, 
                           A1 => n975, B0 => n2759, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831680_127845936_127847840, Y 
                           => n2760);
   U2083 : INVX1 port map( A => n3036, Y => n1054);
   U2084 : AOI22X1 port map( A0 => n1062, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
                           B0 => n3035, B1 => n1055, Y => n3036);
   U2085 : INVX1 port map( A => n2994, Y => n1077);
   U2086 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127715536_127848576, 
                           A1 => n1134, B0 => n2993, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831680_127845936_127847840, Y 
                           => n2994);
   U2087 : INVX1 port map( A => n3504, Y => n577);
   U2088 : AOI22X1 port map( A0 => n585, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
                           B0 => n3503, B1 => n578, Y => n3504);
   U2089 : INVX1 port map( A => n3462, Y => n600);
   U2090 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127715536_127848576, 
                           A1 => n657, B0 => n3461, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831680_127845936_127847840, Y 
                           => n3462);
   U2091 : INVX1 port map( A => n2568, Y => n736);
   U2092 : AOI22X1 port map( A0 => n744, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715648_127848688_127850592, 
                           B0 => n2567, B1 => n737, Y => n2568);
   U2093 : INVX1 port map( A => n2526, Y => n759);
   U2094 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127715536_127848576, 
                           A1 => n816, B0 => n2525, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831680_127845936_127847840, Y 
                           => n2526);
   U2095 : INVX1 port map( A => n4506, Y => n1043);
   U2096 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_15, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_15_port, 
                           B1 => n4495, Y => n4506);
   U2097 : XNOR2X1 port map( A => n3769, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_15, 
                           Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_15_port);
   U2098 : INVX1 port map( A => n4612, Y => n566);
   U2099 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_15,
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_15_port, 
                           B1 => n4601, Y => n4612);
   U2100 : XNOR2X1 port map( A => n3865, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_15,
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_15_port);
   U2101 : INVX1 port map( A => n4505, Y => n1035);
   U2102 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_16, 
                           A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_16_port, 
                           B1 => n4495, Y => n4505);
   U2103 : XNOR2X1 port map( A => n3768, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_16, 
                           Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_16_port);
   U2104 : INVX1 port map( A => n4611, Y => n558);
   U2105 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_16,
                           A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_16_port, 
                           B1 => n4601, Y => n4611);
   U2106 : XNOR2X1 port map( A => n3864, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_16,
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_16_port);
   U2107 : INVX1 port map( A => n4457, Y => n917);
   U2108 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_11, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_11_port, 
                           B1 => n4442, Y => n4457);
   U2109 : XOR2X1 port map( A => n3724, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_11, 
                           Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_11_port);
   U2110 : INVX1 port map( A => input_times_b0_mul_componentxn106, Y => n758);
   U2111 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_11, A1 
                           => n121, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_11_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn106);
   U2112 : XOR2X1 port map( A => n3676, B => 
                           input_times_b0_mul_componentxunsigned_output_11, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_11_port);
   U2113 : BUFX3 port map( A => n254, Y => n144);
   U2114 : BUFX3 port map( A => n282, Y => n132);
   U2115 : INVX1 port map( A => n2724, Y => n974);
   U2116 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127672560_127674464, 
                           A1 => n978, B0 => n2723, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830672_127844928_127846832, Y 
                           => n2724);
   U2117 : INVX1 port map( A => n2958, Y => n1133);
   U2118 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127672560_127674464, 
                           A1 => n1137, B0 => n2957, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830672_127844928_127846832, Y 
                           => n2958);
   U2119 : INVX1 port map( A => n3426, Y => n656);
   U2120 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127672560_127674464, 
                           A1 => n660, B0 => n3425, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830672_127844928_127846832, Y 
                           => n3426);
   U2121 : INVX1 port map( A => n2490, Y => n815);
   U2122 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127672560_127674464, 
                           A1 => n819, B0 => n2489, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830672_127844928_127846832, Y 
                           => n2490);
   U2123 : INVX1 port map( A => n2728, Y => n960);
   U2124 : AOI22X1 port map( A0 => n983, A1 => n964, B0 => n2727, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830896_127845152_127847056, Y 
                           => n2728);
   U2125 : INVX1 port map( A => n2962, Y => n1119);
   U2126 : AOI22X1 port map( A0 => n1142, A1 => n1123, B0 => n2961, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830896_127845152_127847056, Y 
                           => n2962);
   U2127 : INVX1 port map( A => n3430, Y => n642);
   U2128 : AOI22X1 port map( A0 => n665, A1 => n646, B0 => n3429, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830896_127845152_127847056, Y 
                           => n3430);
   U2129 : INVX1 port map( A => n2494, Y => n801);
   U2130 : AOI22X1 port map( A0 => n824, A1 => n805, B0 => n2493, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830896_127845152_127847056, Y 
                           => n2494);
   U2131 : INVX1 port map( A => n2790, Y => n936);
   U2132 : AOI22X1 port map( A0 => n945, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635696_127637600, 
                           B0 => n2789, B1 => n938, Y => n2790);
   U2133 : INVX1 port map( A => n2788, Y => n947);
   U2134 : AOI22X1 port map( A0 => n954, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
                           B0 => n2787, B1 => n948, Y => n2788);
   U2135 : INVX1 port map( A => n3024, Y => n1095);
   U2136 : AOI22X1 port map( A0 => n1104, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635696_127637600, 
                           B0 => n3023, B1 => n1097, Y => n3024);
   U2137 : INVX1 port map( A => n3492, Y => n618);
   U2138 : AOI22X1 port map( A0 => n627, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635696_127637600, 
                           B0 => n3491, B1 => n620, Y => n3492);
   U2139 : INVX1 port map( A => n2556, Y => n777);
   U2140 : AOI22X1 port map( A0 => n786, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635696_127637600, 
                           B0 => n2555, B1 => n779, Y => n2556);
   U2141 : INVX1 port map( A => n2554, Y => n788);
   U2142 : AOI22X1 port map( A0 => n795, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732144_127721824_127723728, 
                           B0 => n2553, B1 => n789, Y => n2554);
   U2143 : INVX1 port map( A => n2976, Y => n1083);
   U2144 : AOI22X1 port map( A0 => n1112, A1 => n1086, B0 => n2975, B1 => n1135
                           , Y => n2976);
   U2145 : INVX1 port map( A => n2990, Y => n1111);
   U2146 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
                           B0 => n2989, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715536_127848576, Y 
                           => n2990);
   U2147 : INVX1 port map( A => n3444, Y => n606);
   U2148 : AOI22X1 port map( A0 => n635, A1 => n609, B0 => n3443, B1 => n658, Y
                           => n3444);
   U2149 : INVX1 port map( A => n3458, Y => n634);
   U2150 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636032_127637936_127713632, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732592_127722272_127724176, 
                           B0 => n3457, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715536_127848576, Y 
                           => n3458);
   U2151 : INVX1 port map( A => n2736, Y => n938);
   U2152 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
                           A1 => n989, B0 => n2735, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673120_127675024_127730240, Y 
                           => n2736);
   U2153 : INVX1 port map( A => n2732, Y => n948);
   U2154 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
                           B0 => n2731, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732032_127721712_127723616, Y 
                           => n2732);
   U2155 : INVX1 port map( A => n2970, Y => n1097);
   U2156 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
                           A1 => n1148, B0 => n2969, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673120_127675024_127730240, Y 
                           => n2970);
   U2157 : INVX1 port map( A => n2966, Y => n1107);
   U2158 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
                           B0 => n2965, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732032_127721712_127723616, Y 
                           => n2966);
   U2159 : INVX1 port map( A => n3438, Y => n620);
   U2160 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
                           A1 => n671, B0 => n3437, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673120_127675024_127730240, Y 
                           => n3438);
   U2161 : INVX1 port map( A => n3434, Y => n630);
   U2162 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
                           B0 => n3433, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732032_127721712_127723616, Y 
                           => n3434);
   U2163 : INVX1 port map( A => n2502, Y => n779);
   U2164 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831120_127845376_127847280, 
                           A1 => n830, B0 => n2501, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673120_127675024_127730240, Y 
                           => n2502);
   U2165 : INVX1 port map( A => n2498, Y => n789);
   U2166 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673008_127674912_127730128, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831008_127845264_127847168, 
                           B0 => n2497, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732032_127721712_127723616, Y 
                           => n2498);
   U2167 : INVX1 port map( A => n2750, Y => n933);
   U2168 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
                           B0 => n2749, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635920_127637824_127713520, Y 
                           => n2750);
   U2169 : INVX1 port map( A => n2754, Y => n896);
   U2170 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
                           A1 => n981, B0 => n2753, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673568_127675472_127730688, Y 
                           => n2754);
   U2171 : INVX1 port map( A => n2984, Y => n1092);
   U2172 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
                           B0 => n2983, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635920_127637824_127713520, Y 
                           => n2984);
   U2173 : INVX1 port map( A => n2988, Y => n1055);
   U2174 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
                           A1 => n1140, B0 => n2987, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673568_127675472_127730688, Y 
                           => n2988);
   U2175 : INVX1 port map( A => n3452, Y => n615);
   U2176 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
                           B0 => n3451, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635920_127637824_127713520, Y 
                           => n3452);
   U2177 : INVX1 port map( A => n3456, Y => n578);
   U2178 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
                           A1 => n663, B0 => n3455, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673568_127675472_127730688, Y 
                           => n3456);
   U2179 : INVX1 port map( A => n2516, Y => n774);
   U2180 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732480_127722160_127724064, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673456_127675360_127730576, 
                           B0 => n2515, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635920_127637824_127713520, Y 
                           => n2516);
   U2181 : INVX1 port map( A => n2520, Y => n737);
   U2182 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831568_127845824_127847728, 
                           A1 => n822, B0 => n2519, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673568_127675472_127730688, Y 
                           => n2520);
   U2183 : INVX1 port map( A => n2780, Y => n973);
   U2184 : AOI22X1 port map( A0 => n979, A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
                           B0 => n2779, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127826576_127826800_127826968, Y 
                           => n2780);
   U2185 : INVX1 port map( A => n3014, Y => n1132);
   U2186 : AOI22X1 port map( A0 => n1138, A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
                           B0 => n3013, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127826576_127826800_127826968, Y 
                           => n3014);
   U2187 : INVX1 port map( A => n3482, Y => n655);
   U2188 : AOI22X1 port map( A0 => n661, A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
                           B0 => n3481, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127826576_127826800_127826968, Y 
                           => n3482);
   U2189 : INVX1 port map( A => n2546, Y => n814);
   U2190 : AOI22X1 port map( A0 => n820, A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672672_127674576_127729792, 
                           B0 => n2545, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer2_127826576_127826800_127826968, Y 
                           => n2546);
   U2191 : BUFX3 port map( A => n254, Y => n143);
   U2192 : BUFX3 port map( A => n282, Y => n131);
   U2193 : BUFX3 port map( A => n255, Y => n141);
   U2194 : BUFX3 port map( A => n256, Y => n139);
   U2195 : BUFX3 port map( A => n255, Y => n142);
   U2196 : BUFX3 port map( A => n256, Y => n140);
   U2197 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_9, 
                           A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_9_port, 
                           B1 => n4442, Y => n4441);
   U2198 : XNOR2X1 port map( A => n3711, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_9, Y
                           => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_9_port);
   U2199 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_9, 
                           A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_9_port, 
                           B1 => n4495, Y => n4494);
   U2200 : XNOR2X1 port map( A => n3759, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_9, Y
                           => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_9_port);
   U2201 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_9, 
                           A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_9_port, 
                           B1 => n4601, Y => n4600);
   U2202 : XNOR2X1 port map( A => n3855, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_9, 
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_9_port);
   U2203 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_9, A1 
                           => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_9_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn90);
   U2204 : XNOR2X1 port map( A => n3663, B => 
                           input_times_b0_mul_componentxunsigned_output_9, Y =>
                           input_times_b0_mul_componentxunsigned_output_inverted_9_port);
   U2205 : INVX1 port map( A => n4497, Y => n1116);
   U2206 : AOI22X1 port map( A0 => n2332, A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_7_port, 
                           B1 => n4495, Y => n4497);
   U2207 : XOR2X1 port map( A => n3761, B => n2332, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_7_port);
   U2208 : INVX1 port map( A => n4603, Y => n639);
   U2209 : AOI22X1 port map( A0 => n2374, A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_7_port, 
                           B1 => n4601, Y => n4603);
   U2210 : XOR2X1 port map( A => n3857, B => n2374, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_7_port);
   U2211 : INVX1 port map( A => n3008, Y => n1033);
   U2212 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
                           B0 => n3007, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636368_127638272_127713968, Y 
                           => n3008);
   U2213 : INVX1 port map( A => n3476, Y => n556);
   U2214 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
                           B0 => n3475, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636368_127638272_127713968, Y 
                           => n3476);
   U2215 : INVX1 port map( A => n2758, Y => n900);
   U2216 : AOI22X1 port map( A0 => n923, A1 => n902, B0 => n2757, B1 => n951, Y
                           => n2758);
   U2217 : INVX1 port map( A => n2992, Y => n1059);
   U2218 : AOI22X1 port map( A0 => n1082, A1 => n1061, B0 => n2991, B1 => n1110
                           , Y => n2992);
   U2219 : INVX1 port map( A => n3460, Y => n582);
   U2220 : AOI22X1 port map( A0 => n605, A1 => n584, B0 => n3459, B1 => n633, Y
                           => n3460);
   U2221 : INVX1 port map( A => n2524, Y => n741);
   U2222 : AOI22X1 port map( A0 => n764, A1 => n743, B0 => n2523, B1 => n792, Y
                           => n2524);
   U2223 : AOI22X1 port map( A0 => n942, A1 => n886, B0 => n2809, B1 => n882, Y
                           => n2810);
   U2224 : AOI22X1 port map( A0 => n1101, A1 => n1045, B0 => n3043, B1 => n1041
                           , Y => n3044);
   U2225 : AOI22X1 port map( A0 => n624, A1 => n568, B0 => n3511, B1 => n564, Y
                           => n3512);
   U2226 : AOI22X1 port map( A0 => n783, A1 => n727, B0 => n2575, B1 => n723, Y
                           => n2576);
   U2227 : XOR2X1 port map( A => n951, B => n2757, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128224392_128224616_128224784);
   U2228 : XOR2X1 port map( A => n1110, B => n2991, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128224392_128224616_128224784);
   U2229 : XOR2X1 port map( A => n633, B => n3459, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128224392_128224616_128224784);
   U2230 : XOR2X1 port map( A => n792, B => n2523, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128224392_128224616_128224784);
   U2231 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673680_127675584_127730800, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732704_127722384_127724288, Y 
                           => n2995);
   U2232 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673680_127675584_127730800, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732704_127722384_127724288, Y 
                           => n3463);
   U2233 : XOR2X1 port map( A => n904, B => n932, Y => n2751);
   U2234 : XOR2X1 port map( A => n1063, B => n1091, Y => n2985);
   U2235 : XOR2X1 port map( A => n586, B => n614, Y => n3453);
   U2236 : XOR2X1 port map( A => n745, B => n773, Y => n2517);
   U2237 : XOR2X1 port map( A => n902, B => n923, Y => n2757);
   U2238 : XOR2X1 port map( A => n1061, B => n1082, Y => n2991);
   U2239 : XOR2X1 port map( A => n584, B => n605, Y => n3459);
   U2240 : XOR2X1 port map( A => n743, B => n764, Y => n2523);
   U2241 : XOR2X1 port map( A => n886, B => n942, Y => n2809);
   U2242 : XOR2X1 port map( A => n1045, B => n1101, Y => n3043);
   U2243 : XOR2X1 port map( A => n568, B => n624, Y => n3511);
   U2244 : XOR2X1 port map( A => n727, B => n783, Y => n2575);
   U2245 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127827752_127827920);
   U2246 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127731920_127721600, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672896_127674800_127730016, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127827752_127827920);
   U2247 : XOR2X1 port map( A => n962, B => n2751, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128223720_128223944_128224168);
   U2248 : XOR2X1 port map( A => n1121, B => n2985, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128223720_128223944_128224168);
   U2249 : XOR2X1 port map( A => n644, B => n3453, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128223720_128223944_128224168);
   U2250 : XOR2X1 port map( A => n803, B => n2517, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128223720_128223944_128224168);
   U2251 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198024_128197968);
   U2252 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198024_128197968);
   U2253 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198024_128197968);
   U2254 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198024_128197968);
   U2255 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830672_127844928_127846832, B 
                           => n2723, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127826576_127826800_127826968);
   U2256 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830672_127844928_127846832, B 
                           => n2957, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127826576_127826800_127826968);
   U2257 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830672_127844928_127846832, B 
                           => n3425, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127826576_127826800_127826968);
   U2258 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830672_127844928_127846832, B 
                           => n2489, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127826576_127826800_127826968);
   U2259 : XOR2X1 port map( A => n976, B => n2741, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128222376_128222600_128222768);
   U2260 : XOR2X1 port map( A => n1135, B => n2975, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128222376_128222600_128222768);
   U2261 : XOR2X1 port map( A => n658, B => n3443, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128222376_128222600_128222768);
   U2262 : XOR2X1 port map( A => n817, B => n2507, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128222376_128222600_128222768);
   U2263 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732816_127722496_127724400, B 
                           => n2767, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197520_128197632_128197800);
   U2264 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732816_127722496_127724400, B 
                           => n2533, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197520_128197632_128197800);
   U2265 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831904_127846160_127848064, B 
                           => n2771, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198080_128198192_128198360);
   U2266 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831904_127846160_127848064, B 
                           => n3005, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198080_128198192_128198360);
   U2267 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831904_127846160_127848064, B 
                           => n3473, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198080_128198192_128198360);
   U2268 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831904_127846160_127848064, B 
                           => n2537, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198080_128198192_128198360);
   U2269 : OR3XL port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_3_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_4_port, C 
                           => n3717, Y => n3715);
   U2270 : OR3XL port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_3_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_4_port, C 
                           => n3765, Y => n3763);
   U2271 : OR3XL port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_3_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_4_port, C 
                           => n3861, Y => n3859);
   U2272 : OR3XL port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_3_port,
                           B => 
                           input_times_b0_mul_componentxUMxfirst_vector_4_port,
                           C => n3669, Y => n3667);
   U2273 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636368_127638272_127713968, B 
                           => n2773, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198472_128198640_128198808);
   U2274 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636368_127638272_127713968, B 
                           => n3007, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198472_128198640_128198808);
   U2275 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636368_127638272_127713968, B 
                           => n3475, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198472_128198640_128198808);
   U2276 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636368_127638272_127713968, B 
                           => n2539, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198472_128198640_128198808);
   U2277 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_128198024_128197968);
   U2278 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_128198024_128197968);
   U2279 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_128198024_128197968);
   U2280 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715760_127848800_127850704, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636256_127638160_127713856, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer2_128198024_128197968);
   U2281 : INVX1 port map( A => n4444, Y => n957);
   U2282 : AOI22X1 port map( A0 => n2311, A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_7_port, 
                           B1 => n4442, Y => n4444);
   U2283 : XOR2X1 port map( A => n3713, B => n2311, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_7_port);
   U2284 : INVX1 port map( A => input_times_b0_mul_componentxn93, Y => n798);
   U2285 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxAdder_finalxn47, A1 
                           => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_7_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn93);
   U2286 : XOR2X1 port map( A => n3665, B => 
                           input_times_b0_mul_componentxUMxAdder_finalxn47, Y 
                           => 
                           input_times_b0_mul_componentxunsigned_output_inverted_7_port);
   U2287 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_127826128_127826296);
   U2288 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_127826128_127826296);
   U2289 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_127826128_127826296);
   U2290 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer2_127826128_127826296);
   U2291 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n987, Y => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer3_128246112_128246336);
   U2292 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n1146, Y => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer3_128246112_128246336);
   U2293 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n669, Y => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer3_128246112_128246336);
   U2294 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n828, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer3_128246112_128246336);
   U2295 : INVX1 port map( A => n4446, Y => n972);
   U2296 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_5_port, 
                           A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_5_port, 
                           B1 => n4442, Y => n4446);
   U2297 : XOR2X1 port map( A => n3715, B => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_5_port, Y 
                           => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_5_port);
   U2298 : INVX1 port map( A => input_times_b0_mul_componentxn95, Y => n813);
   U2299 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxfirst_vector_5_port,
                           A1 => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_5_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn95);
   U2300 : XOR2X1 port map( A => n3667, B => 
                           input_times_b0_mul_componentxUMxfirst_vector_5_port,
                           Y => 
                           input_times_b0_mul_componentxunsigned_output_inverted_5_port);
   U2301 : INVX1 port map( A => n4443, Y => n950);
   U2302 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_8, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_8_port, 
                           B1 => n4442, Y => n4443);
   U2303 : XOR2X1 port map( A => n3712, B => 
                           input_p1_times_b1_mul_componentxunsigned_output_8, Y
                           => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_8_port);
   U2304 : OR2X2 port map( A => n2311, B => n3713, Y => n3712);
   U2305 : INVX1 port map( A => n4496, Y => n1109);
   U2306 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_8, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_8_port, 
                           B1 => n4495, Y => n4496);
   U2307 : XOR2X1 port map( A => n3760, B => 
                           input_p2_times_b2_mul_componentxunsigned_output_8, Y
                           => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_8_port);
   U2308 : OR2X2 port map( A => n2332, B => n3761, Y => n3760);
   U2309 : INVX1 port map( A => n4602, Y => n632);
   U2310 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_8, 
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_8_port, 
                           B1 => n4601, Y => n4602);
   U2311 : XOR2X1 port map( A => n3856, B => 
                           output_p2_times_a2_mul_componentxunsigned_output_8, 
                           Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_8_port);
   U2312 : OR2X2 port map( A => n2374, B => n3857, Y => n3856);
   U2313 : INVX1 port map( A => input_times_b0_mul_componentxn92, Y => n791);
   U2314 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxunsigned_output_8, A1 
                           => n121, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_8_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn92);
   U2315 : XOR2X1 port map( A => n3664, B => 
                           input_times_b0_mul_componentxunsigned_output_8, Y =>
                           input_times_b0_mul_componentxunsigned_output_inverted_8_port);
   U2316 : OR2X2 port map( A => input_times_b0_mul_componentxUMxAdder_finalxn47
                           , B => n3665, Y => n3664);
   U2317 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_128198976_128199144, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198304_128198528_128198696, Y 
                           => n2814);
   U2318 : XOR2X1 port map( A => n922, B => n2775, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198304_128198528_128198696);
   U2319 : AND2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer2_128198976_128199144);
   U2320 : XOR2X1 port map( A => n921, B => n877, Y => n2775);
   U2321 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_128198976_128199144, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198304_128198528_128198696, Y 
                           => n3048);
   U2322 : XOR2X1 port map( A => n1081, B => n3009, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198304_128198528_128198696);
   U2323 : AND2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer2_128198976_128199144);
   U2324 : XOR2X1 port map( A => n1080, B => n1036, Y => n3009);
   U2325 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_128198976_128199144, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198304_128198528_128198696, Y 
                           => n3516);
   U2326 : XOR2X1 port map( A => n604, B => n3477, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198304_128198528_128198696);
   U2327 : AND2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer2_128198976_128199144);
   U2328 : XOR2X1 port map( A => n603, B => n559, Y => n3477);
   U2329 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxcarry_layer2_128198976_128199144, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198304_128198528_128198696, Y 
                           => n2580);
   U2330 : XOR2X1 port map( A => n763, B => n2541, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198304_128198528_128198696);
   U2331 : AND2X2 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer2_128198976_128199144);
   U2332 : XOR2X1 port map( A => n762, B => n718, Y => n2541);
   U2333 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128198976_128199144);
   U2334 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128198976_128199144);
   U2335 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128198976_128199144);
   U2336 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127627504_127629408, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715872_127848912_127850816, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer2_128198976_128199144);
   U2337 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672560_127674464, B 
                           => n2721, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127826464_127826632_127826744);
   U2338 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830448_127844704_127846608, B 
                           => n2719, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127672448_127826240_127826520);
   U2339 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672560_127674464, B 
                           => n2955, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127826464_127826632_127826744);
   U2340 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830448_127844704_127846608, B 
                           => n2953, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127672448_127826240_127826520);
   U2341 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672560_127674464, B 
                           => n3423, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127826464_127826632_127826744);
   U2342 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830448_127844704_127846608, B 
                           => n3421, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127672448_127826240_127826520);
   U2343 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672560_127674464, B 
                           => n2487, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127826464_127826632_127826744);
   U2344 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830448_127844704_127846608, B 
                           => n2485, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_127672448_127826240_127826520);
   U2345 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n987, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer3_128246112_128246336);
   U2346 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n1146, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer3_128246112_128246336);
   U2347 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n669, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer3_128246112_128246336);
   U2348 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer2_127826464_127826632_127826744, B 
                           => n828, Y => 
                           input_times_b0_mul_componentxUMxsum_layer3_128246112_128246336);
   U2349 : INVX1 port map( A => n4445, Y => n965);
   U2350 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_6_port, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_6_port, 
                           B1 => n4442, Y => n4445);
   U2351 : XOR2X1 port map( A => n3714, B => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_6_port, Y 
                           => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_6_port);
   U2352 : OR2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_5_port, B 
                           => n3715, Y => n3714);
   U2353 : INVX1 port map( A => n4498, Y => n1124);
   U2354 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_6_port, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_6_port, 
                           B1 => n4495, Y => n4498);
   U2355 : XOR2X1 port map( A => n3762, B => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_6_port, Y 
                           => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_6_port);
   U2356 : OR2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_5_port, B 
                           => n3763, Y => n3762);
   U2357 : INVX1 port map( A => n4604, Y => n647);
   U2358 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_6_port, 
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_6_port, 
                           B1 => n4601, Y => n4604);
   U2359 : XOR2X1 port map( A => n3858, B => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_6_port, Y 
                           => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_6_port);
   U2360 : OR2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_5_port, B 
                           => n3859, Y => n3858);
   U2361 : INVX1 port map( A => input_times_b0_mul_componentxn94, Y => n806);
   U2362 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxfirst_vector_6_port,
                           A1 => n121, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_6_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn94);
   U2363 : XOR2X1 port map( A => n3666, B => 
                           input_times_b0_mul_componentxUMxfirst_vector_6_port,
                           Y => 
                           input_times_b0_mul_componentxunsigned_output_inverted_6_port);
   U2364 : OR2X2 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_5_port,
                           B => n3667, Y => n3666);
   U2365 : INVX1 port map( A => n2752, Y => n903);
   U2366 : AOI22X1 port map( A0 => n932, A1 => n904, B0 => n2751, B1 => n962, Y
                           => n2752);
   U2367 : INVX1 port map( A => n2986, Y => n1062);
   U2368 : AOI22X1 port map( A0 => n1091, A1 => n1063, B0 => n2985, B1 => n1121
                           , Y => n2986);
   U2369 : INVX1 port map( A => n3454, Y => n585);
   U2370 : AOI22X1 port map( A0 => n614, A1 => n586, B0 => n3453, B1 => n644, Y
                           => n3454);
   U2371 : INVX1 port map( A => n2518, Y => n744);
   U2372 : AOI22X1 port map( A0 => n773, A1 => n745, B0 => n2517, B1 => n803, Y
                           => n2518);
   U2373 : INVX1 port map( A => n2766, Y => n942);
   U2374 : AOI22X1 port map( A0 => n967, A1 => n943, B0 => n2765, B1 => n991, Y
                           => n2766);
   U2375 : INVX1 port map( A => n3000, Y => n1101);
   U2376 : AOI22X1 port map( A0 => n1126, A1 => n1102, B0 => n2999, B1 => n1150
                           , Y => n3000);
   U2377 : INVX1 port map( A => n3468, Y => n624);
   U2378 : AOI22X1 port map( A0 => n649, A1 => n625, B0 => n3467, B1 => n673, Y
                           => n3468);
   U2379 : INVX1 port map( A => n2532, Y => n783);
   U2380 : AOI22X1 port map( A0 => n808, A1 => n784, B0 => n2531, B1 => n832, Y
                           => n2532);
   U2381 : INVX1 port map( A => n2762, Y => n889);
   U2382 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
                           B0 => n2761, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636144_127638048_127713744, Y 
                           => n2762);
   U2383 : INVX1 port map( A => n2996, Y => n1048);
   U2384 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
                           B0 => n2995, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636144_127638048_127713744, Y 
                           => n2996);
   U2385 : INVX1 port map( A => n3464, Y => n571);
   U2386 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
                           B0 => n3463, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636144_127638048_127713744, Y 
                           => n3464);
   U2387 : INVX1 port map( A => n2528, Y => n730);
   U2388 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732704_127722384_127724288, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673680_127675584_127730800, 
                           B0 => n2527, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636144_127638048_127713744, Y 
                           => n2528);
   U2389 : INVX1 port map( A => n2774, Y => n874);
   U2390 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
                           B0 => n2773, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636368_127638272_127713968, Y 
                           => n2774);
   U2391 : INVX1 port map( A => n2540, Y => n715);
   U2392 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732928_127722608_127724512, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673904_127675808_127731024, 
                           B0 => n2539, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636368_127638272_127713968, Y 
                           => n2540);
   U2393 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_2_port);
   U2394 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_2_port);
   U2395 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_2_port);
   U2396 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830336_127844592_127846496, B 
                           => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127830168_127844480, Y 
                           => 
                           input_times_b0_mul_componentxUMxfirst_vector_2_port)
                           ;
   U2397 : XOR2X1 port map( A => n931, B => n2769, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128197464_128197688_128197856);
   U2398 : XOR2X1 port map( A => n1090, B => n3003, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197464_128197688_128197856);
   U2399 : XOR2X1 port map( A => n613, B => n3471, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197464_128197688_128197856);
   U2400 : XOR2X1 port map( A => n772, B => n2535, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128197464_128197688_128197856);
   U2401 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831792_127846048_127847952, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673792_127675696_127730912, Y 
                           => n2767);
   U2402 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831792_127846048_127847952, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673792_127675696_127730912, Y 
                           => n3001);
   U2403 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831792_127846048_127847952, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673792_127675696_127730912, Y 
                           => n3469);
   U2404 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831792_127846048_127847952, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673792_127675696_127730912, Y 
                           => n2533);
   U2405 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673904_127675808_127731024, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732928_127722608_127724512, Y 
                           => n2773);
   U2406 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673904_127675808_127731024, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732928_127722608_127724512, Y 
                           => n3007);
   U2407 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673904_127675808_127731024, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732928_127722608_127724512, Y 
                           => n3475);
   U2408 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673904_127675808_127731024, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732928_127722608_127724512, Y 
                           => n2539);
   U2409 : XOR2X1 port map( A => n920, B => n879, Y => n2769);
   U2410 : XOR2X1 port map( A => n1079, B => n1038, Y => n3003);
   U2411 : XOR2X1 port map( A => n602, B => n561, Y => n3471);
   U2412 : XOR2X1 port map( A => n761, B => n720, Y => n2535);
   U2413 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732816_127722496_127724400, B 
                           => n3001, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128197520_128197632_128197800);
   U2414 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732816_127722496_127724400, B 
                           => n3469, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128197520_128197632_128197800);
   U2415 : OR3XL port map( A => n994, B => n993, C => n995, Y => n3917);
   U2416 : OR3XL port map( A => n1153, B => n1152, C => n1154, Y => n3960);
   U2417 : OR3XL port map( A => n676, B => n675, C => n677, Y => n4046);
   U2418 : OR3XL port map( A => n835, B => n834, C => n836, Y => n3874);
   U2419 : INVX1 port map( A => n4448, Y => n986);
   U2420 : AOI22XL port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_3_port, 
                           A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_3_port, 
                           B1 => n4442, Y => n4448);
   U2421 : XOR2X1 port map( A => n3717, B => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_3_port, Y 
                           => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_3_port);
   U2422 : INVX1 port map( A => n4501, Y => n1145);
   U2423 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_3_port, 
                           A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_3_port, 
                           B1 => n4495, Y => n4501);
   U2424 : XOR2X1 port map( A => n3765, B => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_3_port, Y 
                           => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_3_port);
   U2425 : INVX1 port map( A => n4499, Y => n1131);
   U2426 : AOI22XL port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_5_port, 
                           A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_5_port, 
                           B1 => n4495, Y => n4499);
   U2427 : XOR2X1 port map( A => n3763, B => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_5_port, Y 
                           => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_5_port);
   U2428 : INVX1 port map( A => n4607, Y => n668);
   U2429 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_3_port, 
                           A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_3_port, 
                           B1 => n4601, Y => n4607);
   U2430 : XOR2X1 port map( A => n3861, B => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_3_port, Y 
                           => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_3_port);
   U2431 : INVX1 port map( A => n4605, Y => n654);
   U2432 : AOI22XL port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_5_port, 
                           A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_5_port, 
                           B1 => n4601, Y => n4605);
   U2433 : XOR2X1 port map( A => n3859, B => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_5_port, Y 
                           => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_5_port);
   U2434 : INVX1 port map( A => input_times_b0_mul_componentxn97, Y => n827);
   U2435 : AOI22XL port map( A0 => 
                           input_times_b0_mul_componentxUMxfirst_vector_3_port,
                           A1 => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_3_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn97);
   U2436 : XOR2X1 port map( A => n3669, B => 
                           input_times_b0_mul_componentxUMxfirst_vector_3_port,
                           Y => 
                           input_times_b0_mul_componentxunsigned_output_inverted_3_port);
   U2437 : INVX1 port map( A => n4447, Y => n980);
   U2438 : AOI22XL port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_4_port, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_4_port, 
                           B1 => n4442, Y => n4447);
   U2439 : XOR2X1 port map( A => n3716, B => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_4_port, Y 
                           => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_4_port);
   U2440 : OR2X2 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_3_port, B 
                           => n3717, Y => n3716);
   U2441 : INVX1 port map( A => n4500, Y => n1139);
   U2442 : AOI22XL port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_4_port, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_4_port, 
                           B1 => n4495, Y => n4500);
   U2443 : XOR2X1 port map( A => n3764, B => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_4_port, Y 
                           => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_4_port);
   U2444 : OR2X2 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_3_port, B 
                           => n3765, Y => n3764);
   U2445 : INVX1 port map( A => n4606, Y => n662);
   U2446 : AOI22XL port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_4_port, 
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_4_port, 
                           B1 => n4601, Y => n4606);
   U2447 : XOR2X1 port map( A => n3860, B => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_4_port, Y 
                           => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_4_port);
   U2448 : OR2X2 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_3_port, B 
                           => n3861, Y => n3860);
   U2449 : INVX1 port map( A => input_times_b0_mul_componentxn96, Y => n821);
   U2450 : AOI22XL port map( A0 => 
                           input_times_b0_mul_componentxUMxfirst_vector_4_port,
                           A1 => n121, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_4_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn96);
   U2451 : XOR2X1 port map( A => n3668, B => 
                           input_times_b0_mul_componentxUMxfirst_vector_4_port,
                           Y => 
                           input_times_b0_mul_componentxunsigned_output_inverted_4_port);
   U2452 : OR2X2 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_3_port,
                           B => n3669, Y => n3668);
   U2453 : INVX1 port map( A => n2768, Y => n882);
   U2454 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
                           A1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
                           B0 => n2767, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732816_127722496_127724400, Y 
                           => n2768);
   U2455 : INVX1 port map( A => n3002, Y => n1041);
   U2456 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
                           A1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
                           B0 => n3001, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732816_127722496_127724400, Y 
                           => n3002);
   U2457 : INVX1 port map( A => n3470, Y => n564);
   U2458 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
                           A1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
                           B0 => n3469, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732816_127722496_127724400, Y 
                           => n3470);
   U2459 : INVX1 port map( A => n2534, Y => n723);
   U2460 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673792_127675696_127730912, 
                           A1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831792_127846048_127847952, 
                           B0 => n2533, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732816_127722496_127724400, Y 
                           => n2534);
   U2461 : XNOR2X1 port map( A => n993, B => n3918, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_2_port);
   U2462 : NOR2X1 port map( A => n995, B => n994, Y => n3918);
   U2463 : XNOR2X1 port map( A => n1152, B => n3961, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_2_port);
   U2464 : NOR2X1 port map( A => n1154, B => n1153, Y => n3961);
   U2465 : XNOR2X1 port map( A => n675, B => n4047, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_2_port);
   U2466 : NOR2X1 port map( A => n677, B => n676, Y => n4047);
   U2467 : XNOR2X1 port map( A => n834, B => n3875, Y => 
                           input_times_b0_div_componentxinput_A_inverted_2_port
                           );
   U2468 : NOR2X1 port map( A => n836, B => n835, Y => n3875);
   U2469 : XOR2X1 port map( A => n994, B => n995, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_1_port);
   U2470 : XOR2X1 port map( A => n1153, B => n1154, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_1_port);
   U2471 : XOR2X1 port map( A => n676, B => n677, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_1_port);
   U2472 : XOR2X1 port map( A => n835, B => n836, Y => 
                           input_times_b0_div_componentxinput_A_inverted_1_port
                           );
   U2473 : INVX1 port map( A => n258, Y => n320);
   U2474 : INVX1 port map( A => n258, Y => n319);
   U2475 : INVX1 port map( A => n258, Y => n321);
   U2476 : BUFX3 port map( A => n161, Y => n159);
   U2477 : BUFX3 port map( A => n161, Y => n160);
   U2478 : BUFX3 port map( A => n162, Y => n157);
   U2479 : BUFX3 port map( A => n162, Y => n158);
   U2480 : BUFX3 port map( A => n163, Y => n155);
   U2481 : BUFX3 port map( A => n163, Y => n156);
   U2482 : BUFX3 port map( A => n164, Y => n153);
   U2483 : BUFX3 port map( A => n164, Y => n154);
   U2484 : BUFX3 port map( A => n257, Y => n137);
   U2485 : BUFX3 port map( A => n257, Y => n138);
   U2486 : NOR3X1 port map( A => n853, B => n854, C => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn4, Y 
                           => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn2);
   U2487 : NOR3X1 port map( A => n1012, B => n1013, C => n1762, Y => n1761);
   U2488 : NOR3X1 port map( A => n1171, B => n1172, C => n1771, Y => n1770);
   U2489 : NOR3X1 port map( A => n535, B => n536, C => n1780, Y => n1779);
   U2490 : NOR3X1 port map( A => n694, B => n695, C => n1789, Y => n1788);
   U2491 : NOR3X1 port map( A => output_contracterxn7, B => 
                           output_previous_1_16_port, C => 
                           output_previous_1_15_port, Y => output_contracterxn2
                           );
   U2492 : OR3XL port map( A => n165, B => output_previous_1_8_port, C => 
                           output_previous_1_9_port, Y => output_contracterxn7)
                           ;
   U2493 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn16, B 
                           => n838, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_11_port);
   U2494 : XOR2X1 port map( A => n1768, B => n997, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_11_port);
   U2495 : XOR2X1 port map( A => n1777, B => n1156, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_11_port);
   U2496 : XOR2X1 port map( A => n1786, B => n520, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_11_port);
   U2497 : XOR2X1 port map( A => n1795, B => n679, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_11_port);
   U2498 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn4, B 
                           => n853, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_7_port);
   U2499 : XOR2X1 port map( A => n1762, B => n1012, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_7_port);
   U2500 : XOR2X1 port map( A => n1771, B => n1171, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_7_port);
   U2501 : XOR2X1 port map( A => n1780, B => n535, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_7_port);
   U2502 : XOR2X1 port map( A => n1789, B => n694, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_7_port);
   U2503 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn14, B 
                           => n840, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_13_port);
   U2504 : XOR2X1 port map( A => n1767, B => n999, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_13_port);
   U2505 : XOR2X1 port map( A => n1776, B => n1158, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_13_port);
   U2506 : XOR2X1 port map( A => n1785, B => n522, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_13_port);
   U2507 : XOR2X1 port map( A => n1794, B => n681, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_13_port);
   U2508 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn12, B 
                           => n842, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_15_port);
   U2509 : XOR2X1 port map( A => n1766, B => n1001, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_15_port);
   U2510 : XOR2X1 port map( A => n1775, B => n1160, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_15_port);
   U2511 : XOR2X1 port map( A => n1784, B => n524, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_15_port);
   U2512 : XOR2X1 port map( A => n1793, B => n683, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_15_port);
   U2513 : XNOR2X1 port map( A => n64, B => n854, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_8_port);
   U2514 : NOR2X1 port map( A => n853, B => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn4, Y 
                           => n64);
   U2515 : XNOR2X1 port map( A => n65, B => n1013, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_8_port);
   U2516 : NOR2X1 port map( A => n1012, B => n1762, Y => n65);
   U2517 : XNOR2X1 port map( A => n66, B => n1172, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_8_port);
   U2518 : NOR2X1 port map( A => n1171, B => n1771, Y => n66);
   U2519 : XNOR2X1 port map( A => n67, B => n536, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_8_port);
   U2520 : NOR2X1 port map( A => n535, B => n1780, Y => n67);
   U2521 : XNOR2X1 port map( A => n68, B => n695, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_8_port);
   U2522 : NOR2X1 port map( A => n694, B => n1789, Y => n68);
   U2523 : XNOR2X1 port map( A => n69, B => n839, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_12_port);
   U2524 : NOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn16, B 
                           => n838, Y => n69);
   U2525 : XNOR2X1 port map( A => n70, B => n998, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_12_port);
   U2526 : NOR2X1 port map( A => n1768, B => n997, Y => n70);
   U2527 : XNOR2X1 port map( A => n71, B => n1157, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_12_port);
   U2528 : NOR2X1 port map( A => n1777, B => n1156, Y => n71);
   U2529 : XNOR2X1 port map( A => n72, B => n521, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_12_port);
   U2530 : NOR2X1 port map( A => n1786, B => n520, Y => n72);
   U2531 : XNOR2X1 port map( A => n73, B => n680, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_12_port);
   U2532 : NOR2X1 port map( A => n1795, B => n679, Y => n73);
   U2533 : XNOR2X1 port map( A => n74, B => n841, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_14_port);
   U2534 : NOR2X1 port map( A => n840, B => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn14, Y 
                           => n74);
   U2535 : XNOR2X1 port map( A => n75, B => n1000, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_14_port);
   U2536 : NOR2X1 port map( A => n999, B => n1767, Y => n75);
   U2537 : XNOR2X1 port map( A => n76, B => n1159, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_14_port);
   U2538 : NOR2X1 port map( A => n1158, B => n1776, Y => n76);
   U2539 : XNOR2X1 port map( A => n77, B => n523, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_14_port);
   U2540 : NOR2X1 port map( A => n522, B => n1785, Y => n77);
   U2541 : XNOR2X1 port map( A => n78, B => n682, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_14_port);
   U2542 : NOR2X1 port map( A => n681, B => n1794, Y => n78);
   U2543 : OR3XL port map( A => n838, B => n839, C => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn16, Y 
                           => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn14);
   U2544 : OR3XL port map( A => n997, B => n998, C => n1768, Y => n1767);
   U2545 : OR3XL port map( A => n1156, B => n1157, C => n1777, Y => n1776);
   U2546 : OR3XL port map( A => n520, B => n521, C => n1786, Y => n1785);
   U2547 : OR3XL port map( A => n679, B => n680, C => n1795, Y => n1794);
   U2548 : NAND3X1 port map( A => output_previous_1_16_port, B => 
                           output_previous_1_15_port, C => n165, Y => 
                           output_contracterxn6);
   U2549 : OR3XL port map( A => n840, B => n841, C => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn14, Y 
                           => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn12);
   U2550 : OR3XL port map( A => n999, B => n1000, C => n1767, Y => n1766);
   U2551 : OR3XL port map( A => n1158, B => n1159, C => n1776, Y => n1775);
   U2552 : OR3XL port map( A => n522, B => n523, C => n1785, Y => n1784);
   U2553 : OR3XL port map( A => n681, B => n682, C => n1794, Y => n1793);
   U2554 : BUFX3 port map( A => output_previous_1_17_port, Y => n165);
   U2555 : XOR2X1 port map( A => n4169, B => n4170, Y => 
                           output_previous_1_17_port);
   U2556 : XNOR2X1 port map( A => results_a1_a2_inv_17_port, B => 
                           results_b0_b1_b2_17_port, Y => n4169);
   U2557 : AOI22X1 port map( A0 => n4171, A1 => n1205, B0 => 
                           results_b0_b1_b2_16_port, B1 => 
                           results_a1_a2_inv_16_port, Y => n4170);
   U2558 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b4,
                           B => output_p1_times_a1_mul_componentxUMxa1_and_b3, 
                           Y => n3095);
   U2559 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b5,
                           B => output_p1_times_a1_mul_componentxUMxa1_and_b4, 
                           Y => n3097);
   U2560 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b0,
                           B => n494, Y => n3193);
   U2561 : XOR2X1 port map( A => n4121, B => n4122, Y => results_a1_a2_8_port);
   U2562 : XOR2X1 port map( A => results_b0_b1_adderxn14, B => 
                           results_b0_b1_adderxn15, Y => results_b0_b1_3_port);
   U2563 : XOR2X1 port map( A => n4098, B => n4099, Y => 
                           results_b0_b1_b2_3_port);
   U2564 : XOR2X1 port map( A => results_b0_b1_adderxn10, B => 
                           results_b0_b1_adderxn11, Y => results_b0_b1_5_port);
   U2565 : XOR2X1 port map( A => n4094, B => n4095, Y => 
                           results_b0_b1_b2_5_port);
   U2566 : XOR2X1 port map( A => results_b0_b1_adderxn6, B => 
                           results_b0_b1_adderxn7, Y => results_b0_b1_7_port);
   U2567 : XOR2X1 port map( A => n4090, B => n4091, Y => 
                           results_b0_b1_b2_7_port);
   U2568 : XOR2X1 port map( A => results_b0_b1_adderxn2, B => 
                           results_b0_b1_adderxn3, Y => results_b0_b1_9_port);
   U2569 : XOR2X1 port map( A => n4086, B => n4087, Y => 
                           results_b0_b1_b2_9_port);
   U2570 : XOR2X1 port map( A => results_b0_b1_adderxn32, B => 
                           results_b0_b1_adderxn33, Y => results_b0_b1_11_port)
                           ;
   U2571 : XOR2X1 port map( A => n4115, B => n4116, Y => 
                           results_b0_b1_b2_11_port);
   U2572 : XOR2X1 port map( A => results_b0_b1_adderxn28, B => 
                           results_b0_b1_adderxn29, Y => results_b0_b1_13_port)
                           ;
   U2573 : XOR2X1 port map( A => n4111, B => n4112, Y => 
                           results_b0_b1_b2_13_port);
   U2574 : XOR2X1 port map( A => n4107, B => n4108, Y => 
                           results_b0_b1_b2_15_port);
   U2575 : XOR2X1 port map( A => n4125, B => n4126, Y => results_a1_a2_6_port);
   U2576 : XOR2X1 port map( A => results_b0_b1_adderxn16, B => 
                           results_b0_b1_adderxn17, Y => results_b0_b1_2_port);
   U2577 : XOR2X1 port map( A => n4100, B => n4101, Y => 
                           results_b0_b1_b2_2_port);
   U2578 : XOR2X1 port map( A => results_b0_b1_adderxn12, B => 
                           results_b0_b1_adderxn13, Y => results_b0_b1_4_port);
   U2579 : XOR2X1 port map( A => n4096, B => n4097, Y => 
                           results_b0_b1_b2_4_port);
   U2580 : XOR2X1 port map( A => results_b0_b1_adderxn8, B => 
                           results_b0_b1_adderxn9, Y => results_b0_b1_6_port);
   U2581 : XOR2X1 port map( A => n4092, B => n4093, Y => 
                           results_b0_b1_b2_6_port);
   U2582 : XOR2X1 port map( A => results_b0_b1_adderxn4, B => 
                           results_b0_b1_adderxn5, Y => results_b0_b1_8_port);
   U2583 : XOR2X1 port map( A => n4088, B => n4089, Y => 
                           results_b0_b1_b2_8_port);
   U2584 : XOR2X1 port map( A => results_b0_b1_adderxn35, B => 
                           results_b0_b1_adderxn34, Y => results_b0_b1_10_port)
                           ;
   U2585 : XOR2X1 port map( A => n4118, B => n4117, Y => 
                           results_b0_b1_b2_10_port);
   U2586 : XOR2X1 port map( A => results_b0_b1_adderxn31, B => 
                           results_b0_b1_adderxn30, Y => results_b0_b1_12_port)
                           ;
   U2587 : XOR2X1 port map( A => n4114, B => n4113, Y => 
                           results_b0_b1_b2_12_port);
   U2588 : XOR2X1 port map( A => results_b0_b1_adderxn27, B => 
                           results_b0_b1_adderxn26, Y => results_b0_b1_14_port)
                           ;
   U2589 : XOR2X1 port map( A => n4110, B => n4109, Y => 
                           results_b0_b1_b2_14_port);
   U2590 : INVX1 port map( A => n3098, Y => n494);
   U2591 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b4, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b5, B0 =>
                           n3097, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b3, Y => 
                           n3098);
   U2592 : INVX1 port map( A => n3096, Y => n501);
   U2593 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b3, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b4, B0 =>
                           n3095, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b2, Y => 
                           n3096);
   U2594 : INVX1 port map( A => n3194, Y => n493);
   U2595 : AOI22X1 port map( A0 => n494, A1 => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b0, B0 =>
                           n3193, B1 => n513, Y => n3194);
   U2596 : BUFX3 port map( A => n1321, Y => n146);
   U2597 : BUFX3 port map( A => n1341, Y => n148);
   U2598 : BUFX3 port map( A => n1380, Y => n152);
   U2599 : BUFX3 port map( A => n1238, Y => n136);
   U2600 : AOI32X1 port map( A0 => results_a1_a2_inv_0_port, A1 => n4168, A2 =>
                           results_b0_b1_b2_0_port, B0 => 
                           results_a1_a2_inv_1_port, B1 => 
                           results_b0_b1_b2_1_port, Y => n4167);
   U2601 : NOR2X1 port map( A => n4528, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b10);
   U2602 : NOR2X1 port map( A => n4527, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b11);
   U2603 : NOR2X1 port map( A => n4526, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b12);
   U2604 : NOR2X1 port map( A => n214, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b7);
   U2605 : NOR2X1 port map( A => n213, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b8);
   U2606 : NOR2X1 port map( A => n212, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b9);
   U2607 : NOR2X1 port map( A => n213, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b8);
   U2608 : NOR2X1 port map( A => n214, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b7);
   U2609 : INVX1 port map( A => n3142, Y => n504);
   U2610 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b2, A1 
                           => output_p1_times_a1_mul_componentxUMxa9_and_b3, B0
                           => n3141, B1 => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b1, Y =>
                           n3142);
   U2611 : NOR2X1 port map( A => n231, B => n4528, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b10);
   U2612 : NOR2X1 port map( A => n231, B => n4527, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b11);
   U2613 : INVX1 port map( A => n3094, Y => n508);
   U2614 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b2, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b3, B0 =>
                           n3093, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b1, Y => 
                           n3094);
   U2615 : INVX1 port map( A => n3108, Y => n500);
   U2616 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b3, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b4, B0 =>
                           n3107, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b2, Y => 
                           n3108);
   U2617 : INVX1 port map( A => n3106, Y => n479);
   U2618 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b6, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b7, B0 =>
                           n3105, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b5, Y => 
                           n3106);
   U2619 : INVX1 port map( A => n3092, Y => n515);
   U2620 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b1, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b2, B0 =>
                           n3091, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b0, Y => 
                           n3092);
   U2621 : INVX1 port map( A => n3102, Y => n487);
   U2622 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b5, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b6, B0 =>
                           n3101, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b4, Y => 
                           n3102);
   U2623 : INVX1 port map( A => n3110, Y => n469);
   U2624 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b7, A1 =>
                           output_p1_times_a1_mul_componentxUMxa0_and_b8, B0 =>
                           n3109, B1 => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b6, Y => 
                           n3110);
   U2625 : INVX1 port map( A => n3114, Y => n512);
   U2626 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b1, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b2, B0 =>
                           n3113, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b0, Y => 
                           n3114);
   U2627 : INVX1 port map( A => n3132, Y => n491);
   U2628 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b4, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b5, B0 =>
                           n3131, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b3, Y => 
                           n3132);
   U2629 : NOR2X1 port map( A => n231, B => n4526, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b12);
   U2630 : NOR2X1 port map( A => n231, B => n4525, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b13);
   U2631 : NOR2X1 port map( A => n231, B => n214, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b7);
   U2632 : NOR2X1 port map( A => n231, B => n213, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b8);
   U2633 : NOR2X1 port map( A => n231, B => n212, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b9);
   U2634 : NOR2X1 port map( A => n212, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b9);
   U2635 : NOR2X1 port map( A => n214, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b7);
   U2636 : NOR2X1 port map( A => n214, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b7);
   U2637 : NOR2X1 port map( A => n213, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b8);
   U2638 : XOR2X1 port map( A => n4123, B => n4124, Y => results_a1_a2_7_port);
   U2639 : XOR2X1 port map( A => n4144, B => n4145, Y => results_a1_a2_13_port)
                           ;
   U2640 : XOR2X1 port map( A => n4119, B => n4120, Y => results_a1_a2_9_port);
   U2641 : XOR2X1 port map( A => n4131, B => n4132, Y => results_a1_a2_3_port);
   U2642 : XOR2X1 port map( A => n4127, B => n4128, Y => results_a1_a2_5_port);
   U2643 : XOR2X1 port map( A => n4148, B => n4149, Y => results_a1_a2_11_port)
                           ;
   U2644 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b2,
                           B => n3095, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830560_127844816_127846720);
   U2645 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b3,
                           B => n3111, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673008_127674912_127730128);
   U2646 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b4,
                           B => n3139, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732480_127722160_127724064);
   U2647 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b5,
                           B => n3123, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673232_127675136_127730352);
   U2648 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa12_and_b0
                           , B => n436, Y => n3213);
   U2649 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b3,
                           B => output_p1_times_a1_mul_componentxUMxa1_and_b2, 
                           Y => n3093);
   U2650 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b7,
                           B => output_p1_times_a1_mul_componentxUMxa1_and_b6, 
                           Y => n3105);
   U2651 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b2,
                           B => output_p1_times_a1_mul_componentxUMxa1_and_b1, 
                           Y => n3091);
   U2652 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b6,
                           B => output_p1_times_a1_mul_componentxUMxa1_and_b5, 
                           Y => n3101);
   U2653 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b0,
                           B => n515, Y => n3187);
   U2654 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa9_and_b0,
                           B => n469, Y => n3201);
   U2655 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b2,
                           B => output_p1_times_a1_mul_componentxUMxa4_and_b1, 
                           Y => n3099);
   U2656 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b2,
                           B => output_p1_times_a1_mul_componentxUMxa7_and_b1, 
                           Y => n3113);
   U2657 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b3,
                           B => output_p1_times_a1_mul_componentxUMxa4_and_b2, 
                           Y => n3103);
   U2658 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b3,
                           B => output_p1_times_a1_mul_componentxUMxa7_and_b2, 
                           Y => n3119);
   U2659 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b4,
                           B => output_p1_times_a1_mul_componentxUMxa4_and_b3, 
                           Y => n3107);
   U2660 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b4,
                           B => output_p1_times_a1_mul_componentxUMxa7_and_b3, 
                           Y => n3125);
   U2661 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b5,
                           B => output_p1_times_a1_mul_componentxUMxa4_and_b4, 
                           Y => n3111);
   U2662 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b5,
                           B => output_p1_times_a1_mul_componentxUMxa7_and_b4, 
                           Y => n3131);
   U2663 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa9_and_b2,
                           B => output_p1_times_a1_mul_componentxUMxa10_and_b1,
                           Y => n3133);
   U2664 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa9_and_b3,
                           B => output_p1_times_a1_mul_componentxUMxa10_and_b2,
                           Y => n3141);
   U2665 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b6,
                           B => output_p1_times_a1_mul_componentxUMxa4_and_b5, 
                           Y => n3117);
   U2666 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b7,
                           B => output_p1_times_a1_mul_componentxUMxa4_and_b6, 
                           Y => n3123);
   U2667 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b6,
                           B => output_p1_times_a1_mul_componentxUMxa7_and_b5, 
                           Y => n3139);
   U2668 : XOR2X1 port map( A => n4140, B => n4141, Y => results_a1_a2_15_port)
                           ;
   U2669 : XOR2X1 port map( A => n4143, B => n4142, Y => results_a1_a2_14_port)
                           ;
   U2670 : AND2X2 port map( A => output_p1_times_a1_mul_componentxUMxa4_and_b0,
                           B => output_p1_times_a1_mul_componentxUMxa3_and_b1, 
                           Y => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127672560_127674464);
   U2671 : XOR2X1 port map( A => results_b0_b1_b2_1_port, B => 
                           results_a1_a2_inv_1_port, Y => n4168);
   U2672 : XOR2X1 port map( A => results_a1_a2_1_port, B => 
                           results_a1_a2_inv_0_port, Y => 
                           results_a1_a2_inv_1_port);
   U2673 : XNOR2X1 port map( A => results_a1_a2_2_port, B => 
                           results_a1_a2_inv_inverterxn9, Y => 
                           results_a1_a2_inv_2_port);
   U2674 : NOR2X1 port map( A => results_a1_a2_inv_0_port, B => 
                           results_a1_a2_1_port, Y => 
                           results_a1_a2_inv_inverterxn9);
   U2675 : XOR2X1 port map( A => results_b0_b1_adderxn24, B => 
                           results_b0_b1_adderxn25, Y => results_b0_b1_15_port)
                           ;
   U2676 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b0,
                           B => n3099, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672672_127674576_127729792);
   U2677 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b1,
                           B => n3119, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732144_127721824_127723728);
   U2678 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b6,
                           B => n3109, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127831008_127845264_127847168);
   U2679 : OR3XL port map( A => results_a1_a2_1_port, B => results_a1_a2_2_port
                           , C => results_a1_a2_inv_0_port, Y => 
                           results_a1_a2_inv_inverterxn8);
   U2680 : XOR2X1 port map( A => n4129, B => n4130, Y => results_a1_a2_4_port);
   U2681 : XOR2X1 port map( A => n4147, B => n4146, Y => results_a1_a2_12_port)
                           ;
   U2682 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b0,
                           B => n3113, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732032_127721712_127723616);
   U2683 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b2,
                           B => n3125, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732256_127721936_127723840);
   U2684 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b3,
                           B => n3097, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830672_127844928_127846832);
   U2685 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b4,
                           B => n3117, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673120_127675024_127730240);
   U2686 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b5,
                           B => n3105, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830896_127845152_127847056);
   U2687 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa4_and_b0,
                           B => output_p1_times_a1_mul_componentxUMxa3_and_b1, 
                           Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672560_127674464);
   U2688 : XOR2X1 port map( A => results_b0_b1_adderxn22, B => n1209, Y => 
                           results_b0_b1_16_port);
   U2689 : XOR2X1 port map( A => n4105, B => n1207, Y => 
                           results_b0_b1_b2_16_port);
   U2690 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b2,
                           B => n3107, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672896_127674800_127730016);
   U2691 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b4,
                           B => n3101, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830784_127845040_127846944);
   U2692 : XOR2X1 port map( A => n4151, B => n4150, Y => results_a1_a2_10_port)
                           ;
   U2693 : XOR2X1 port map( A => n4138, B => n1301, Y => results_a1_a2_16_port)
                           ;
   U2694 : AND2X2 port map( A => output_p1_times_a1_mul_componentxUMxa7_and_b0,
                           B => output_p1_times_a1_mul_componentxUMxa6_and_b1, 
                           Y => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127731920_127721600);
   U2695 : XOR2X1 port map( A => n4133, B => n4134, Y => results_a1_a2_2_port);
   U2696 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b1,
                           B => n3103, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127672784_127674688_127729904);
   U2697 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa7_and_b0,
                           B => output_p1_times_a1_mul_componentxUMxa6_and_b1, 
                           Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127731920_127721600);
   U2698 : INVX1 port map( A => n3134, Y => n511);
   U2699 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b1, A1 
                           => output_p1_times_a1_mul_componentxUMxa9_and_b2, B0
                           => n3133, B1 => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b0, Y =>
                           n3134);
   U2700 : INVX1 port map( A => n3104, Y => n506);
   U2701 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b2, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b3, B0 =>
                           n3103, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b1, Y => 
                           n3104);
   U2702 : INVX1 port map( A => n3118, Y => n486);
   U2703 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b5, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b6, B0 =>
                           n3117, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b4, Y => 
                           n3118);
   U2704 : INVX1 port map( A => n3202, Y => n468);
   U2705 : AOI22X1 port map( A0 => n469, A1 => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b0, B0 =>
                           n3201, B1 => n492, Y => n3202);
   U2706 : INVX1 port map( A => n3124, Y => n476);
   U2707 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b6, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b7, B0 =>
                           n3123, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b5, Y => 
                           n3124);
   U2708 : BUFX3 port map( A => n1321, Y => n145);
   U2709 : BUFX3 port map( A => n1341, Y => n147);
   U2710 : BUFX3 port map( A => n1380, Y => n151);
   U2711 : BUFX3 port map( A => n1238, Y => n135);
   U2712 : BUFX3 port map( A => n1360, Y => n149);
   U2713 : INVX1 port map( A => n3214, Y => n435);
   U2714 : AOI22X1 port map( A0 => n436, A1 => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b0, B0 
                           => n3213, B1 => n467, Y => n3214);
   U2715 : INVX1 port map( A => n3100, Y => n513);
   U2716 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b1, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b2, B0 =>
                           n3099, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b0, Y => 
                           n3100);
   U2717 : INVX1 port map( A => n3112, Y => n492);
   U2718 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b4, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b5, B0 =>
                           n3111, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b3, Y => 
                           n3112);
   U2719 : INVX1 port map( A => n3130, Y => n467);
   U2720 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b7, A1 =>
                           output_p1_times_a1_mul_componentxUMxa3_and_b8, B0 =>
                           n3129, B1 => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b6, Y => 
                           n3130);
   U2721 : INVX1 port map( A => n3120, Y => n505);
   U2722 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b2, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b3, B0 =>
                           n3119, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b1, Y => 
                           n3120);
   U2723 : INVX1 port map( A => n3188, Y => n510);
   U2724 : AOI22X1 port map( A0 => n515, A1 => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b0, B0 =>
                           n3187, B1 => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830448_127844704_127846608, Y 
                           => n3188);
   U2725 : BUFX3 port map( A => n1360, Y => n150);
   U2726 : NAND2X1 port map( A => results_b0_b1_b2_0_port, B => 
                           results_a1_a2_inv_0_port, Y => n79);
   U2727 : NOR2X1 port map( A => n4528, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b10);
   U2728 : NOR2X1 port map( A => n4527, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b11);
   U2729 : NOR2X1 port map( A => n4525, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b13);
   U2730 : NOR2X1 port map( A => n4524, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b14);
   U2731 : NOR2X1 port map( A => n212, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b9);
   U2732 : NOR2X1 port map( A => n214, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b7);
   U2733 : NOR2X1 port map( A => n4528, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b10);
   U2734 : INVX1 port map( A => n3150, Y => n498);
   U2735 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b3, A1 
                           => output_p1_times_a1_mul_componentxUMxa9_and_b4, B0
                           => n3149, B1 => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b2, Y =>
                           n3150);
   U2736 : NOR2X1 port map( A => n4528, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b10);
   U2737 : NOR2X1 port map( A => n4527, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b11);
   U2738 : NOR2X1 port map( A => n4527, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b11);
   U2739 : NOR2X1 port map( A => n4526, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b12);
   U2740 : NOR2X1 port map( A => n4526, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b12);
   U2741 : NOR2X1 port map( A => n231, B => n4524, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b14);
   U2742 : NOR2X1 port map( A => n231, B => n4523, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b15);
   U2743 : NOR2X1 port map( A => n213, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b8);
   U2744 : NOR2X1 port map( A => n214, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b7);
   U2745 : NOR2X1 port map( A => n213, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b8);
   U2746 : NOR2X1 port map( A => n212, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b9);
   U2747 : NOR2X1 port map( A => n214, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b7);
   U2748 : NOR2X1 port map( A => n213, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b8);
   U2749 : NOR2X1 port map( A => n212, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b9);
   U2750 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa11_and_b2
                           , B => n3149, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636032_127637936_127713632);
   U2751 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b6,
                           B => n3155, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732704_127722384_127724288);
   U2752 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa12_and_b2
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b1, Y =>
                           n3159);
   U2753 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa12_and_b3
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b2, Y =>
                           n3169);
   U2754 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa15_and_b0
                           , B => n443, Y => n3231);
   U2755 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa9_and_b4,
                           B => output_p1_times_a1_mul_componentxUMxa10_and_b3,
                           Y => n3149);
   U2756 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b7,
                           B => output_p1_times_a1_mul_componentxUMxa7_and_b6, 
                           Y => n3147);
   U2757 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa9_and_b5,
                           B => output_p1_times_a1_mul_componentxUMxa10_and_b4,
                           Y => n3157);
   U2758 : AND2X2 port map( A => output_p1_times_a1_mul_componentxUMxa13_and_b0
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b1, Y =>
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127715536_127848576);
   U2759 : OR3XL port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_1_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_2_port, C 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_0_port, Y 
                           => n3813);
   U2760 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa14_and_b0
                           , B => n3159, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715648_127848688_127850592);
   U2761 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b5,
                           B => n3147, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732592_127722272_127724176);
   U2762 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa10_and_b0
                           , B => output_p1_times_a1_mul_componentxUMxa9_and_b1
                           , Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635696_127637600);
   U2763 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa11_and_b1
                           , B => n3141, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635920_127637824_127713520);
   U2764 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa11_and_b3
                           , B => n3157, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636144_127638048_127713744);
   U2765 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b1,
                           B => n3093, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830448_127844704_127846608);
   U2766 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b6,
                           B => n3129, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127673344_127675248_127730464);
   U2767 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa13_and_b0
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b1, Y =>
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715536_127848576);
   U2768 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b3,
                           B => n3131, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127732368_127722048_127723952);
   U2769 : AND2X2 port map( A => output_p1_times_a1_mul_componentxUMxa10_and_b0
                           , B => output_p1_times_a1_mul_componentxUMxa9_and_b1
                           , Y => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127635696_127637600);
   U2770 : AND2X2 port map( A => output_p1_times_a1_mul_componentxUMxa1_and_b0,
                           B => output_p1_times_a1_mul_componentxUMxa0_and_b1, 
                           Y => 
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127830168_127844480);
   U2771 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa11_and_b0
                           , B => n3133, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127635808_127637712_127713408);
   U2772 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b0,
                           B => n3091, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127830336_127844592_127846496);
   U2773 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128238312_128238424_128238592, B 
                           => n405, Y => n3324);
   U2774 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128264344_128264512, B 
                           => n3304, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer4_128238312_128238424_128238592);
   U2775 : INVX1 port map( A => n3318, Y => n405);
   U2776 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128199816_128200040_128199984, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128199368_128199480_128199648, Y 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer3_128264344_128264512);
   U2777 : INVX1 port map( A => n3158, Y => n490);
   U2778 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b4, A1 
                           => output_p1_times_a1_mul_componentxUMxa9_and_b5, B0
                           => n3157, B1 => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b3, Y =>
                           n3158);
   U2779 : INVX1 port map( A => n3170, Y => n507);
   U2780 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b2, A1 
                           => output_p1_times_a1_mul_componentxUMxa12_and_b3, 
                           B0 => n3169, B1 => 
                           output_p1_times_a1_mul_componentxUMxa14_and_b1, Y =>
                           n3170);
   U2781 : INVX1 port map( A => n3156, Y => n466);
   U2782 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b7, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b8, B0 =>
                           n3155, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b6, Y => 
                           n3156);
   U2783 : INVX1 port map( A => n3160, Y => n514);
   U2784 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b1, A1 
                           => output_p1_times_a1_mul_componentxUMxa12_and_b2, 
                           B0 => n3159, B1 => 
                           output_p1_times_a1_mul_componentxUMxa14_and_b0, Y =>
                           n3160);
   U2785 : INVX1 port map( A => n3140, Y => n485);
   U2786 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b5, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b6, B0 =>
                           n3139, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b4, Y => 
                           n3140);
   U2787 : INVX1 port map( A => n3126, Y => n499);
   U2788 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b3, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b4, B0 =>
                           n3125, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b2, Y => 
                           n3126);
   U2789 : INVX1 port map( A => n3148, Y => n474);
   U2790 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b6, A1 =>
                           output_p1_times_a1_mul_componentxUMxa6_and_b7, B0 =>
                           n3147, B1 => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b5, Y => 
                           n3148);
   U2791 : NOR2X1 port map( A => n4526, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b12);
   U2792 : NOR2X1 port map( A => n4523, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b15);
   U2793 : NOR2X1 port map( A => n213, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b8);
   U2794 : NOR2X1 port map( A => n212, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b9);
   U2795 : NOR2X1 port map( A => n4528, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b10);
   U2796 : INVX1 port map( A => n3168, Y => n484);
   U2797 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b5, A1 
                           => output_p1_times_a1_mul_componentxUMxa9_and_b6, B0
                           => n3167, B1 => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b4, Y =>
                           n3168);
   U2798 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b3, A1 
                           => output_p1_times_a1_mul_componentxUMxa12_and_b4, 
                           B0 => n3179, B1 => 
                           output_p1_times_a1_mul_componentxUMxa14_and_b2, Y =>
                           n3180);
   U2799 : NOR2X1 port map( A => n4528, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b10);
   U2800 : NOR2X1 port map( A => n4527, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b11);
   U2801 : NOR2X1 port map( A => n4525, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b13);
   U2802 : NOR2X1 port map( A => n4525, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b13);
   U2803 : NOR2X1 port map( A => n4524, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b14);
   U2804 : NOR2X1 port map( A => n231, B => n4522, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b16);
   U2805 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa1_and_b0,
                           B => output_p1_times_a1_mul_componentxUMxa0_and_b1, 
                           Y => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_1_port);
   U2806 : NOR2X1 port map( A => n212, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b9);
   U2807 : NOR2X1 port map( A => n222, B => n214, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b7);
   U2808 : NOR2X1 port map( A => n214, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b7);
   U2809 : NOR2X1 port map( A => n213, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b8);
   U2810 : NOR2X1 port map( A => n214, B => n4545, Y => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b7);
   U2811 : NOR2X1 port map( A => n4525, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b13);
   U2812 : NOR2X1 port map( A => n4522, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b16);
   U2813 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa12_and_b4
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b3, Y =>
                           n3179);
   U2814 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa9_and_b6,
                           B => output_p1_times_a1_mul_componentxUMxa10_and_b5,
                           Y => n3167);
   U2815 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa9_and_b7,
                           B => output_p1_times_a1_mul_componentxUMxa10_and_b6,
                           Y => n3177);
   U2816 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa11_and_b5
                           , B => n3177, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636368_127638272_127713968);
   U2817 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa11_and_b4
                           , B => n3167, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636256_127638160_127713856);
   U2818 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa14_and_b2
                           , B => n3179, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715872_127848912_127850816);
   U2819 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa14_and_b1
                           , B => n3169, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715760_127848800_127850704);
   U2820 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa16_and_b0
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa15_and_b1, Y =>
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127627504_127629408);
   U2821 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa5_and_b12
                           , B => n3182, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127674016_127675920_127731136);
   U2822 : NOR2X1 port map( A => n4526, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b12);
   U2823 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa3_and_b14
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b13, Y =>
                           n3182);
   U2824 : NOR2X1 port map( A => n4524, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b14);
   U2825 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127733040_127722720_127724624, B 
                           => n3245, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128199368_128199480_128199648);
   U2826 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa8_and_b9,
                           B => n3183, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127733040_127722720_127724624);
   U2827 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127832016_127846272_127848176, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127674016_127675920_127731136, Y 
                           => n3245);
   U2828 : NOR2X1 port map( A => n212, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b9);
   U2829 : XOR2X1 port map( A => n3178, B => n3180, Y => n3244);
   U2830 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b6, A1 
                           => output_p1_times_a1_mul_componentxUMxa9_and_b7, B0
                           => n3177, B1 => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b5, Y =>
                           n3178);
   U2831 : INVX1 port map( A => n4555, Y => n516);
   U2832 : AOI22XL port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_2_port, 
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_2_port, 
                           B1 => n4548, Y => n4555);
   U2833 : XNOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_2_port, B 
                           => n3814, Y => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_2_port);
   U2834 : NOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_0_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_1_port, Y 
                           => n3814);
   U2835 : INVX1 port map( A => n4556, Y => n517);
   U2836 : AOI22XL port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_1_port, 
                           A1 => n114, B0 => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_1_port, 
                           B1 => n4548, Y => n4556);
   U2837 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_1_port, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_0_port, Y 
                           => 
                           output_p1_times_a1_mul_componentxunsigned_output_inverted_1_port);
   U2838 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa2_and_b15
                           , B => n3181, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127832016_127846272_127848176);
   U2839 : NOR2X1 port map( A => n4523, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b15);
   U2840 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa0_and_b17
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b16, Y =>
                           n3181);
   U2841 : NOR2X1 port map( A => n231, B => n20, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b17);
   U2842 : INVX1 port map( A => n3232, Y => n410);
   U2843 : AOI22X1 port map( A0 => n443, A1 => 
                           output_p1_times_a1_mul_componentxUMxa15_and_b0, B0 
                           => n3231, B1 => n411, Y => n3232);
   U2844 : AND2X2 port map( A => output_p1_times_a1_mul_componentxUMxa16_and_b0
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa15_and_b1, Y =>
                           output_p1_times_a1_mul_componentxUMxcarry_layer1_127627504_127629408);
   U2845 : INVX1 port map( A => n4565, Y => n518);
   U2846 : AOI22XL port map( A0 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_0_port, 
                           A1 => n113, B0 => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_0_port, 
                           B1 => n4548, Y => n4565);
   U2847 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa6_and_b11
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b10, Y =>
                           n3183);
   U2848 : NOR2X1 port map( A => n4527, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b11);
   U2849 : NOR2X1 port map( A => n4528, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b10);
   U2850 : XOR2X1 port map( A => n134, B => n361, Y => n80);
   U2851 : INVX1 port map( A => n80, Y => n4548);
   U2852 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa9_and_b2, 
                           B => input_p1_times_b1_mul_componentxUMxa10_and_b1, 
                           Y => n2665);
   U2853 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa9_and_b2, 
                           B => input_p2_times_b2_mul_componentxUMxa10_and_b1, 
                           Y => n2899);
   U2854 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa9_and_b2,
                           B => output_p2_times_a2_mul_componentxUMxa10_and_b1,
                           Y => n3367);
   U2855 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa9_and_b2, B 
                           => input_times_b0_mul_componentxUMxa10_and_b1, Y => 
                           n2431);
   U2856 : INVX1 port map( A => n2666, Y => n988);
   U2857 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b1, A1 =>
                           input_p1_times_b1_mul_componentxUMxa9_and_b2, B0 => 
                           n2665, B1 => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b0, Y => 
                           n2666);
   U2858 : INVX1 port map( A => n2900, Y => n1147);
   U2859 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b1, A1 =>
                           input_p2_times_b2_mul_componentxUMxa9_and_b2, B0 => 
                           n2899, B1 => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b0, Y => 
                           n2900);
   U2860 : INVX1 port map( A => n3368, Y => n670);
   U2861 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b1, A1 
                           => output_p2_times_a2_mul_componentxUMxa9_and_b2, B0
                           => n3367, B1 => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b0, Y =>
                           n3368);
   U2862 : INVX1 port map( A => n2432, Y => n829);
   U2863 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa10_and_b1, 
                           A1 => input_times_b0_mul_componentxUMxa9_and_b2, B0 
                           => n2431, B1 => 
                           input_times_b0_mul_componentxUMxa11_and_b0, Y => 
                           n2432);
   U2864 : INVX1 port map( A => n2674, Y => n981);
   U2865 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b2, A1 =>
                           input_p1_times_b1_mul_componentxUMxa9_and_b3, B0 => 
                           n2673, B1 => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b1, Y => 
                           n2674);
   U2866 : INVX1 port map( A => n2440, Y => n822);
   U2867 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa10_and_b2, 
                           A1 => input_times_b0_mul_componentxUMxa9_and_b3, B0 
                           => n2439, B1 => 
                           input_times_b0_mul_componentxUMxa11_and_b1, Y => 
                           n2440);
   U2868 : INVX1 port map( A => n2682, Y => n975);
   U2869 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b3, A1 =>
                           input_p1_times_b1_mul_componentxUMxa9_and_b4, B0 => 
                           n2681, B1 => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b2, Y => 
                           n2682);
   U2870 : INVX1 port map( A => n2448, Y => n816);
   U2871 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa10_and_b3, 
                           A1 => input_times_b0_mul_componentxUMxa9_and_b4, B0 
                           => n2447, B1 => 
                           input_times_b0_mul_componentxUMxa11_and_b2, Y => 
                           n2448);
   U2872 : INVX1 port map( A => n2628, Y => n978);
   U2873 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b3
                           , A1 => input_p1_times_b1_mul_componentxUMxa0_and_b4
                           , B0 => n2627, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b2, Y => 
                           n2628);
   U2874 : INVX1 port map( A => n2862, Y => n1137);
   U2875 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b3
                           , A1 => input_p2_times_b2_mul_componentxUMxa0_and_b4
                           , B0 => n2861, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b2, Y => 
                           n2862);
   U2876 : INVX1 port map( A => n3330, Y => n660);
   U2877 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b3, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b4, B0 =>
                           n3329, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b2, Y => 
                           n3330);
   U2878 : INVX1 port map( A => n2394, Y => n819);
   U2879 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b3, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b4, B0 
                           => n2393, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b2, Y => 
                           n2394);
   U2880 : INVX1 port map( A => n2630, Y => n971);
   U2881 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b4
                           , A1 => input_p1_times_b1_mul_componentxUMxa0_and_b5
                           , B0 => n2629, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b3, Y => 
                           n2630);
   U2882 : INVX1 port map( A => n2396, Y => n812);
   U2883 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b4, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b5, B0 
                           => n2395, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b3, Y => 
                           n2396);
   U2884 : INVX1 port map( A => n2860, Y => n1144);
   U2885 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b2
                           , A1 => input_p2_times_b2_mul_componentxUMxa0_and_b3
                           , B0 => n2859, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b1, Y => 
                           n2860);
   U2886 : INVX1 port map( A => n3328, Y => n667);
   U2887 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b2, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b3, B0 =>
                           n3327, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b1, Y => 
                           n3328);
   U2888 : INVX1 port map( A => n2636, Y => n983);
   U2889 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b2
                           , A1 => input_p1_times_b1_mul_componentxUMxa3_and_b3
                           , B0 => n2635, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b1, Y => 
                           n2636);
   U2890 : INVX1 port map( A => n2874, Y => n1136);
   U2891 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b3
                           , A1 => input_p2_times_b2_mul_componentxUMxa3_and_b4
                           , B0 => n2873, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b2, Y => 
                           n2874);
   U2892 : INVX1 port map( A => n2872, Y => n1115);
   U2893 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b6
                           , A1 => input_p2_times_b2_mul_componentxUMxa0_and_b7
                           , B0 => n2871, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b5, Y => 
                           n2872);
   U2894 : INVX1 port map( A => n3342, Y => n659);
   U2895 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b3, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b4, B0 =>
                           n3341, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b2, Y => 
                           n3342);
   U2896 : INVX1 port map( A => n3340, Y => n638);
   U2897 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b6, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b7, B0 =>
                           n3339, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b5, Y => 
                           n3340);
   U2898 : INVX1 port map( A => n2402, Y => n824);
   U2899 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b2, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b3, B0 
                           => n2401, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b1, Y => 
                           n2402);
   U2900 : INVX1 port map( A => n2726, Y => n970);
   U2901 : AOI22X1 port map( A0 => n971, A1 => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b0, B0 => 
                           n2725, B1 => n990, Y => n2726);
   U2902 : INVX1 port map( A => n2646, Y => n989);
   U2903 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b1
                           , A1 => input_p1_times_b1_mul_componentxUMxa6_and_b2
                           , B0 => n2645, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b0, Y => 
                           n2646);
   U2904 : INVX1 port map( A => n2960, Y => n1129);
   U2905 : AOI22X1 port map( A0 => n1130, A1 => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b0, B0 => 
                           n2959, B1 => n1149, Y => n2960);
   U2906 : INVX1 port map( A => n3428, Y => n652);
   U2907 : AOI22X1 port map( A0 => n653, A1 => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b0, B0 =>
                           n3427, B1 => n672, Y => n3428);
   U2908 : INVX1 port map( A => n2492, Y => n811);
   U2909 : AOI22X1 port map( A0 => n812, A1 => 
                           input_times_b0_mul_componentxUMxa6_and_b0, B0 => 
                           n2491, B1 => n831, Y => n2492);
   U2910 : INVX1 port map( A => n2412, Y => n830);
   U2911 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b1, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b2, B0 
                           => n2411, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b0, Y => 
                           n2412);
   U2912 : INVX1 port map( A => n2734, Y => n945);
   U2913 : AOI22X1 port map( A0 => n946, A1 => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b0, B0 => 
                           n2733, B1 => n969, Y => n2734);
   U2914 : INVX1 port map( A => n2664, Y => n968);
   U2915 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b4
                           , A1 => input_p1_times_b1_mul_componentxUMxa6_and_b5
                           , B0 => n2663, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b3, Y => 
                           n2664);
   U2916 : INVX1 port map( A => n2898, Y => n1127);
   U2917 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b4
                           , A1 => input_p2_times_b2_mul_componentxUMxa6_and_b5
                           , B0 => n2897, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b3, Y => 
                           n2898);
   U2918 : INVX1 port map( A => n3366, Y => n650);
   U2919 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b4, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b5, B0 =>
                           n3365, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b3, Y => 
                           n3366);
   U2920 : INVX1 port map( A => n2500, Y => n786);
   U2921 : AOI22X1 port map( A0 => n787, A1 => 
                           input_times_b0_mul_componentxUMxa9_and_b0, B0 => 
                           n2499, B1 => n810, Y => n2500);
   U2922 : INVX1 port map( A => n2430, Y => n809);
   U2923 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b4, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b5, B0 
                           => n2429, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b3, Y => 
                           n2430);
   U2924 : INVX1 port map( A => n2656, Y => n953);
   U2925 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b6
                           , A1 => input_p1_times_b1_mul_componentxUMxa3_and_b7
                           , B0 => n2655, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b5, Y => 
                           n2656);
   U2926 : INVX1 port map( A => n2422, Y => n794);
   U2927 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b6, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b7, B0 
                           => n2421, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b5, Y => 
                           n2422);
   U2928 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa11_and_b2,
                           B => n2681, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636032_127637936_127713632);
   U2929 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa11_and_b2, B 
                           => n2447, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636032_127637936_127713632);
   U2930 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa11_and_b2,
                           B => n2915, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636032_127637936_127713632);
   U2931 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa11_and_b2
                           , B => n3383, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636032_127637936_127713632);
   U2932 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b2, 
                           B => n2627, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830560_127844816_127846720);
   U2933 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b2, 
                           B => n2861, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830560_127844816_127846720);
   U2934 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b2,
                           B => n3329, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830560_127844816_127846720);
   U2935 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b2, B 
                           => n2393, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830560_127844816_127846720);
   U2936 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b3, 
                           B => n2643, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673008_127674912_127730128);
   U2937 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b3, 
                           B => n2877, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673008_127674912_127730128);
   U2938 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b3,
                           B => n3345, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673008_127674912_127730128);
   U2939 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b3, B 
                           => n2409, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673008_127674912_127730128);
   U2940 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b4, 
                           B => n2671, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732480_127722160_127724064);
   U2941 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b4, 
                           B => n2905, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732480_127722160_127724064);
   U2942 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b4,
                           B => n3373, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732480_127722160_127724064);
   U2943 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b4, B 
                           => n2437, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732480_127722160_127724064);
   U2944 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b5, 
                           B => n2655, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673232_127675136_127730352);
   U2945 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b5, 
                           B => n2889, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673232_127675136_127730352);
   U2946 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b5,
                           B => n3357, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673232_127675136_127730352);
   U2947 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b5, B 
                           => n2421, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673232_127675136_127730352);
   U2948 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b6, 
                           B => n2687, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732704_127722384_127724288);
   U2949 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b6, B 
                           => n2453, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732704_127722384_127724288);
   U2950 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa12_and_b0,
                           B => n912, Y => n2745);
   U2951 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa12_and_b0, B 
                           => n753, Y => n2511);
   U2952 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa12_and_b2,
                           B => input_p1_times_b1_mul_componentxUMxa13_and_b1, 
                           Y => n2691);
   U2953 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa12_and_b2, B 
                           => input_times_b0_mul_componentxUMxa13_and_b1, Y => 
                           n2457);
   U2954 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa12_and_b3,
                           B => input_p1_times_b1_mul_componentxUMxa13_and_b2, 
                           Y => n2701);
   U2955 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa12_and_b3, B 
                           => input_times_b0_mul_componentxUMxa13_and_b2, Y => 
                           n2467);
   U2956 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa12_and_b0,
                           B => n1071, Y => n2979);
   U2957 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa12_and_b0
                           , B => n594, Y => n3447);
   U2958 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa12_and_b2,
                           B => input_p2_times_b2_mul_componentxUMxa13_and_b1, 
                           Y => n2925);
   U2959 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa12_and_b2
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b1, Y =>
                           n3393);
   U2960 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa12_and_b3,
                           B => input_p2_times_b2_mul_componentxUMxa13_and_b2, 
                           Y => n2935);
   U2961 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa12_and_b3
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b2, Y =>
                           n3403);
   U2962 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa15_and_b0,
                           B => n919, Y => n2763);
   U2963 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa15_and_b0, B 
                           => n760, Y => n2529);
   U2964 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa15_and_b0,
                           B => n1078, Y => n2997);
   U2965 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa15_and_b0
                           , B => n601, Y => n3465);
   U2966 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b4, 
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b3, Y
                           => n2627);
   U2967 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b4, 
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b3, Y
                           => n2861);
   U2968 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b4,
                           B => output_p2_times_a2_mul_componentxUMxa1_and_b3, 
                           Y => n3329);
   U2969 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b4, B 
                           => input_times_b0_mul_componentxUMxa1_and_b3, Y => 
                           n2393);
   U2970 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b5, 
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b4, Y
                           => n2629);
   U2971 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b5, 
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b4, Y
                           => n2863);
   U2972 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b5,
                           B => output_p2_times_a2_mul_componentxUMxa1_and_b4, 
                           Y => n3331);
   U2973 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b5, B 
                           => input_times_b0_mul_componentxUMxa1_and_b4, Y => 
                           n2395);
   U2974 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b3, 
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b2, Y
                           => n2625);
   U2975 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b3, 
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b2, Y
                           => n2859);
   U2976 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b3,
                           B => output_p2_times_a2_mul_componentxUMxa1_and_b2, 
                           Y => n3327);
   U2977 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b3, B 
                           => input_times_b0_mul_componentxUMxa1_and_b2, Y => 
                           n2391);
   U2978 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b8, 
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b7, Y
                           => n2641);
   U2979 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b7, 
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b6, Y
                           => n2637);
   U2980 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b8, 
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b7, Y
                           => n2875);
   U2981 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b7, 
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b6, Y
                           => n2871);
   U2982 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b8,
                           B => output_p2_times_a2_mul_componentxUMxa1_and_b7, 
                           Y => n3343);
   U2983 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b7,
                           B => output_p2_times_a2_mul_componentxUMxa1_and_b6, 
                           Y => n3339);
   U2984 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b8, B 
                           => input_times_b0_mul_componentxUMxa1_and_b7, Y => 
                           n2407);
   U2985 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b7, B 
                           => input_times_b0_mul_componentxUMxa1_and_b6, Y => 
                           n2403);
   U2986 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b0, 
                           B => n971, Y => n2725);
   U2987 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b6, 
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b5, Y
                           => n2633);
   U2988 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b0, 
                           B => n1130, Y => n2959);
   U2989 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b6, 
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b5, Y
                           => n2867);
   U2990 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b0,
                           B => n653, Y => n3427);
   U2991 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b6,
                           B => output_p2_times_a2_mul_componentxUMxa1_and_b5, 
                           Y => n3335);
   U2992 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b0, B 
                           => n812, Y => n2491);
   U2993 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b6, B 
                           => input_times_b0_mul_componentxUMxa1_and_b5, Y => 
                           n2399);
   U2994 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa9_and_b0, 
                           B => n946, Y => n2733);
   U2995 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa9_and_b0, 
                           B => n1105, Y => n2967);
   U2996 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa9_and_b0,
                           B => n628, Y => n3435);
   U2997 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa9_and_b0, B 
                           => n787, Y => n2499);
   U2998 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b2, 
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b1, Y
                           => n2631);
   U2999 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b2, 
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b1, Y
                           => n2865);
   U3000 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b2,
                           B => output_p2_times_a2_mul_componentxUMxa4_and_b1, 
                           Y => n3333);
   U3001 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b2, B 
                           => input_times_b0_mul_componentxUMxa4_and_b1, Y => 
                           n2397);
   U3002 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b2, 
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b1, Y
                           => n2645);
   U3003 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b2, 
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b1, Y
                           => n2879);
   U3004 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b2,
                           B => output_p2_times_a2_mul_componentxUMxa7_and_b1, 
                           Y => n3347);
   U3005 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b2, B 
                           => input_times_b0_mul_componentxUMxa7_and_b1, Y => 
                           n2411);
   U3006 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b3, 
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b2, Y
                           => n2635);
   U3007 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b3, 
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b2, Y
                           => n2869);
   U3008 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b3,
                           B => output_p2_times_a2_mul_componentxUMxa4_and_b2, 
                           Y => n3337);
   U3009 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b3, B 
                           => input_times_b0_mul_componentxUMxa4_and_b2, Y => 
                           n2401);
   U3010 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b3, 
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b2, Y
                           => n2651);
   U3011 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b3, 
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b2, Y
                           => n2885);
   U3012 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b3,
                           B => output_p2_times_a2_mul_componentxUMxa7_and_b2, 
                           Y => n3353);
   U3013 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b3, B 
                           => input_times_b0_mul_componentxUMxa7_and_b2, Y => 
                           n2417);
   U3014 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b4, 
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b3, Y
                           => n2639);
   U3015 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b4, 
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b3, Y
                           => n2873);
   U3016 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b4,
                           B => output_p2_times_a2_mul_componentxUMxa4_and_b3, 
                           Y => n3341);
   U3017 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b4, B 
                           => input_times_b0_mul_componentxUMxa4_and_b3, Y => 
                           n2405);
   U3018 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b4, 
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b3, Y
                           => n2657);
   U3019 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b4, 
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b3, Y
                           => n2891);
   U3020 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b4,
                           B => output_p2_times_a2_mul_componentxUMxa7_and_b3, 
                           Y => n3359);
   U3021 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b4, B 
                           => input_times_b0_mul_componentxUMxa7_and_b3, Y => 
                           n2423);
   U3022 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b5, 
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b4, Y
                           => n2643);
   U3023 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b5, 
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b4, Y
                           => n2877);
   U3024 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b5,
                           B => output_p2_times_a2_mul_componentxUMxa4_and_b4, 
                           Y => n3345);
   U3025 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b5, B 
                           => input_times_b0_mul_componentxUMxa4_and_b4, Y => 
                           n2409);
   U3026 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b5, 
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b4, Y
                           => n2663);
   U3027 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b5, 
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b4, Y
                           => n2897);
   U3028 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b5,
                           B => output_p2_times_a2_mul_componentxUMxa7_and_b4, 
                           Y => n3365);
   U3029 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b5, B 
                           => input_times_b0_mul_componentxUMxa7_and_b4, Y => 
                           n2429);
   U3030 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b6, 
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b5, Y
                           => n2649);
   U3031 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b6, 
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b5, Y
                           => n2883);
   U3032 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b6,
                           B => output_p2_times_a2_mul_componentxUMxa4_and_b5, 
                           Y => n3351);
   U3033 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b6, B 
                           => input_times_b0_mul_componentxUMxa4_and_b5, Y => 
                           n2415);
   U3034 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b6, 
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b5, Y
                           => n2671);
   U3035 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b6, 
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b5, Y
                           => n2905);
   U3036 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b6,
                           B => output_p2_times_a2_mul_componentxUMxa7_and_b5, 
                           Y => n3373);
   U3037 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b6, B 
                           => input_times_b0_mul_componentxUMxa7_and_b5, Y => 
                           n2437);
   U3038 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b7, 
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b6, Y
                           => n2655);
   U3039 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa9_and_b3, 
                           B => input_p1_times_b1_mul_componentxUMxa10_and_b2, 
                           Y => n2673);
   U3040 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b7, 
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b6, Y
                           => n2889);
   U3041 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa9_and_b3, 
                           B => input_p2_times_b2_mul_componentxUMxa10_and_b2, 
                           Y => n2907);
   U3042 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b7,
                           B => output_p2_times_a2_mul_componentxUMxa4_and_b6, 
                           Y => n3357);
   U3043 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa9_and_b3,
                           B => output_p2_times_a2_mul_componentxUMxa10_and_b2,
                           Y => n3375);
   U3044 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b7, B 
                           => input_times_b0_mul_componentxUMxa4_and_b6, Y => 
                           n2421);
   U3045 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa9_and_b3, B 
                           => input_times_b0_mul_componentxUMxa10_and_b2, Y => 
                           n2439);
   U3046 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa9_and_b4, 
                           B => input_p1_times_b1_mul_componentxUMxa10_and_b3, 
                           Y => n2681);
   U3047 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa9_and_b4, 
                           B => input_p2_times_b2_mul_componentxUMxa10_and_b3, 
                           Y => n2915);
   U3048 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa9_and_b4,
                           B => output_p2_times_a2_mul_componentxUMxa10_and_b3,
                           Y => n3383);
   U3049 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa9_and_b4, B 
                           => input_times_b0_mul_componentxUMxa10_and_b3, Y => 
                           n2447);
   U3050 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa9_and_b5, 
                           B => input_p1_times_b1_mul_componentxUMxa10_and_b4, 
                           Y => n2689);
   U3051 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa9_and_b5, 
                           B => input_p2_times_b2_mul_componentxUMxa10_and_b4, 
                           Y => n2923);
   U3052 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa9_and_b5,
                           B => output_p2_times_a2_mul_componentxUMxa10_and_b4,
                           Y => n3391);
   U3053 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa9_and_b5, B 
                           => input_times_b0_mul_componentxUMxa10_and_b4, Y => 
                           n2455);
   U3054 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b8, 
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b7, Y
                           => n2687);
   U3055 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b8, B 
                           => input_times_b0_mul_componentxUMxa7_and_b7, Y => 
                           n2453);
   U3056 : AND2X2 port map( A => input_p1_times_b1_mul_componentxUMxa13_and_b0,
                           B => input_p1_times_b1_mul_componentxUMxa12_and_b1, 
                           Y => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127715536_127848576);
   U3057 : AND2X2 port map( A => input_times_b0_mul_componentxUMxa13_and_b0, B 
                           => input_times_b0_mul_componentxUMxa12_and_b1, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127715536_127848576);
   U3058 : AND2X2 port map( A => input_p2_times_b2_mul_componentxUMxa13_and_b0,
                           B => input_p2_times_b2_mul_componentxUMxa12_and_b1, 
                           Y => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127715536_127848576);
   U3059 : AND2X2 port map( A => output_p2_times_a2_mul_componentxUMxa13_and_b0
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b1, Y =>
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127715536_127848576);
   U3060 : AND2X2 port map( A => input_p1_times_b1_mul_componentxUMxa4_and_b0, 
                           B => input_p1_times_b1_mul_componentxUMxa3_and_b1, Y
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127672560_127674464);
   U3061 : AND2X2 port map( A => input_p2_times_b2_mul_componentxUMxa4_and_b0, 
                           B => input_p2_times_b2_mul_componentxUMxa3_and_b1, Y
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127672560_127674464);
   U3062 : AND2X2 port map( A => output_p2_times_a2_mul_componentxUMxa4_and_b0,
                           B => output_p2_times_a2_mul_componentxUMxa3_and_b1, 
                           Y => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127672560_127674464);
   U3063 : AND2X2 port map( A => input_times_b0_mul_componentxUMxa4_and_b0, B 
                           => input_times_b0_mul_componentxUMxa3_and_b1, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127672560_127674464);
   U3064 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa14_and_b0,
                           B => n2691, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715648_127848688_127850592);
   U3065 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa14_and_b0, B 
                           => n2457, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715648_127848688_127850592);
   U3066 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa14_and_b0,
                           B => n2925, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715648_127848688_127850592);
   U3067 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa14_and_b0
                           , B => n3393, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715648_127848688_127850592);
   U3068 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b1, 
                           B => n2651, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732144_127721824_127723728);
   U3069 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b1, 
                           B => n2885, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732144_127721824_127723728);
   U3070 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b1,
                           B => n3353, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732144_127721824_127723728);
   U3071 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b1, B 
                           => n2417, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732144_127721824_127723728);
   U3072 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b6, 
                           B => n2641, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831008_127845264_127847168);
   U3073 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b6, 
                           B => n2875, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831008_127845264_127847168);
   U3074 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b6,
                           B => n3343, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831008_127845264_127847168);
   U3075 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b6, B 
                           => n2407, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831008_127845264_127847168);
   U3076 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa10_and_b0,
                           B => input_p1_times_b1_mul_componentxUMxa9_and_b1, Y
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635696_127637600);
   U3077 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa10_and_b0,
                           B => input_p2_times_b2_mul_componentxUMxa9_and_b1, Y
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635696_127637600);
   U3078 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa10_and_b0
                           , B => output_p2_times_a2_mul_componentxUMxa9_and_b1
                           , Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635696_127637600);
   U3079 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa10_and_b0, B 
                           => input_times_b0_mul_componentxUMxa9_and_b1, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635696_127637600);
   U3080 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa11_and_b1,
                           B => n2673, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635920_127637824_127713520);
   U3081 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa11_and_b1, B 
                           => n2439, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635920_127637824_127713520);
   U3082 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa11_and_b3,
                           B => n2689, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636144_127638048_127713744);
   U3083 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa11_and_b3, B 
                           => n2455, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636144_127638048_127713744);
   U3084 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa11_and_b1,
                           B => n2907, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635920_127637824_127713520);
   U3085 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa11_and_b1
                           , B => n3375, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635920_127637824_127713520);
   U3086 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa11_and_b3,
                           B => n2923, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636144_127638048_127713744);
   U3087 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa11_and_b3
                           , B => n3391, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636144_127638048_127713744);
   U3088 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b0, 
                           B => n2645, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732032_127721712_127723616);
   U3089 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b0, 
                           B => n2879, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732032_127721712_127723616);
   U3090 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b0,
                           B => n3347, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732032_127721712_127723616);
   U3091 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b0, B 
                           => n2411, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732032_127721712_127723616);
   U3092 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b2, 
                           B => n2657, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732256_127721936_127723840);
   U3093 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b2, 
                           B => n2891, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732256_127721936_127723840);
   U3094 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b2,
                           B => n3359, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732256_127721936_127723840);
   U3095 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b2, B 
                           => n2423, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732256_127721936_127723840);
   U3096 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b3, 
                           B => n2629, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830672_127844928_127846832);
   U3097 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b3, 
                           B => n2863, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830672_127844928_127846832);
   U3098 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b3,
                           B => n3331, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830672_127844928_127846832);
   U3099 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b3, B 
                           => n2395, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830672_127844928_127846832);
   U3100 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b4, 
                           B => n2649, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673120_127675024_127730240);
   U3101 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b4, B 
                           => n2415, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673120_127675024_127730240);
   U3102 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b5, 
                           B => n2637, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830896_127845152_127847056);
   U3103 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b5, 
                           B => n2871, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830896_127845152_127847056);
   U3104 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b5,
                           B => n3339, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830896_127845152_127847056);
   U3105 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b5, B 
                           => n2403, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830896_127845152_127847056);
   U3106 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa13_and_b0,
                           B => input_p1_times_b1_mul_componentxUMxa12_and_b1, 
                           Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715536_127848576);
   U3107 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa13_and_b0, B 
                           => input_times_b0_mul_componentxUMxa12_and_b1, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715536_127848576);
   U3108 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa13_and_b0,
                           B => input_p2_times_b2_mul_componentxUMxa12_and_b1, 
                           Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715536_127848576);
   U3109 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa13_and_b0
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b1, Y =>
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715536_127848576);
   U3110 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b2, 
                           B => n2639, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672896_127674800_127730016);
   U3111 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b2, 
                           B => n2873, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672896_127674800_127730016);
   U3112 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b2,
                           B => n3341, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672896_127674800_127730016);
   U3113 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b2, B 
                           => n2405, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672896_127674800_127730016);
   U3114 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b4, 
                           B => n2633, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830784_127845040_127846944);
   U3115 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b4, 
                           B => n2867, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830784_127845040_127846944);
   U3116 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b4,
                           B => n3335, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830784_127845040_127846944);
   U3117 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b4, B 
                           => n2399, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830784_127845040_127846944);
   U3118 : AND2X2 port map( A => input_p1_times_b1_mul_componentxUMxa10_and_b0,
                           B => input_p1_times_b1_mul_componentxUMxa9_and_b1, Y
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127635696_127637600);
   U3119 : AND2X2 port map( A => input_p2_times_b2_mul_componentxUMxa10_and_b0,
                           B => input_p2_times_b2_mul_componentxUMxa9_and_b1, Y
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127635696_127637600);
   U3120 : AND2X2 port map( A => output_p2_times_a2_mul_componentxUMxa10_and_b0
                           , B => output_p2_times_a2_mul_componentxUMxa9_and_b1
                           , Y => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127635696_127637600);
   U3121 : AND2X2 port map( A => input_times_b0_mul_componentxUMxa10_and_b0, B 
                           => input_times_b0_mul_componentxUMxa9_and_b1, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127635696_127637600);
   U3122 : AND2X2 port map( A => input_p1_times_b1_mul_componentxUMxa7_and_b0, 
                           B => input_p1_times_b1_mul_componentxUMxa6_and_b1, Y
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127731920_127721600);
   U3123 : AND2X2 port map( A => input_p2_times_b2_mul_componentxUMxa7_and_b0, 
                           B => input_p2_times_b2_mul_componentxUMxa6_and_b1, Y
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127731920_127721600);
   U3124 : AND2X2 port map( A => output_p2_times_a2_mul_componentxUMxa7_and_b0,
                           B => output_p2_times_a2_mul_componentxUMxa6_and_b1, 
                           Y => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127731920_127721600);
   U3125 : AND2X2 port map( A => input_times_b0_mul_componentxUMxa7_and_b0, B 
                           => input_times_b0_mul_componentxUMxa6_and_b1, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127731920_127721600);
   U3126 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa11_and_b0,
                           B => n2665, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127635808_127637712_127713408);
   U3127 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa11_and_b0, B 
                           => n2431, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127635808_127637712_127713408);
   U3128 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa11_and_b0,
                           B => n2899, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127635808_127637712_127713408);
   U3129 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa11_and_b0
                           , B => n3367, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127635808_127637712_127713408);
   U3130 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b1, 
                           B => n2635, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672784_127674688_127729904);
   U3131 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b1, 
                           B => n2869, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672784_127674688_127729904);
   U3132 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b1,
                           B => n3337, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672784_127674688_127729904);
   U3133 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b1, B 
                           => n2401, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672784_127674688_127729904);
   U3134 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa7_and_b0, 
                           B => input_p1_times_b1_mul_componentxUMxa6_and_b1, Y
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127731920_127721600);
   U3135 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa7_and_b0, 
                           B => input_p2_times_b2_mul_componentxUMxa6_and_b1, Y
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127731920_127721600);
   U3136 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa7_and_b0,
                           B => output_p2_times_a2_mul_componentxUMxa6_and_b1, 
                           Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127731920_127721600);
   U3137 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa7_and_b0, B 
                           => input_times_b0_mul_componentxUMxa6_and_b1, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127731920_127721600);
   U3138 : INVX1 port map( A => n2690, Y => n967);
   U3139 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b4, A1 =>
                           input_p1_times_b1_mul_componentxUMxa9_and_b5, B0 => 
                           n2689, B1 => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b3, Y => 
                           n2690);
   U3140 : INVX1 port map( A => n2924, Y => n1126);
   U3141 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b4, A1 =>
                           input_p2_times_b2_mul_componentxUMxa9_and_b5, B0 => 
                           n2923, B1 => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b3, Y => 
                           n2924);
   U3142 : INVX1 port map( A => n3392, Y => n649);
   U3143 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b4, A1 
                           => output_p2_times_a2_mul_componentxUMxa9_and_b5, B0
                           => n3391, B1 => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b3, Y =>
                           n3392);
   U3144 : INVX1 port map( A => n2456, Y => n808);
   U3145 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa10_and_b4, 
                           A1 => input_times_b0_mul_componentxUMxa9_and_b5, B0 
                           => n2455, B1 => 
                           input_times_b0_mul_componentxUMxa11_and_b3, Y => 
                           n2456);
   U3146 : INVX1 port map( A => n2702, Y => n984);
   U3147 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa13_and_b2, A1 =>
                           input_p1_times_b1_mul_componentxUMxa12_and_b3, B0 =>
                           n2701, B1 => 
                           input_p1_times_b1_mul_componentxUMxa14_and_b1, Y => 
                           n2702);
   U3148 : INVX1 port map( A => n2936, Y => n1143);
   U3149 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa13_and_b2, A1 =>
                           input_p2_times_b2_mul_componentxUMxa12_and_b3, B0 =>
                           n2935, B1 => 
                           input_p2_times_b2_mul_componentxUMxa14_and_b1, Y => 
                           n2936);
   U3150 : INVX1 port map( A => n3404, Y => n666);
   U3151 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b2, A1 
                           => output_p2_times_a2_mul_componentxUMxa12_and_b3, 
                           B0 => n3403, B1 => 
                           output_p2_times_a2_mul_componentxUMxa14_and_b1, Y =>
                           n3404);
   U3152 : INVX1 port map( A => n2468, Y => n825);
   U3153 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa13_and_b2, 
                           A1 => input_times_b0_mul_componentxUMxa12_and_b3, B0
                           => n2467, B1 => 
                           input_times_b0_mul_componentxUMxa14_and_b1, Y => 
                           n2468);
   U3154 : INVX1 port map( A => n2864, Y => n1130);
   U3155 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b4
                           , A1 => input_p2_times_b2_mul_componentxUMxa0_and_b5
                           , B0 => n2863, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b3, Y => 
                           n2864);
   U3156 : INVX1 port map( A => n3332, Y => n653);
   U3157 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b4, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b5, B0 =>
                           n3331, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b3, Y => 
                           n3332);
   U3158 : INVX1 port map( A => n2642, Y => n946);
   U3159 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b7
                           , A1 => input_p1_times_b1_mul_componentxUMxa0_and_b8
                           , B0 => n2641, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b6, Y => 
                           n2642);
   U3160 : INVX1 port map( A => n2640, Y => n977);
   U3161 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b3
                           , A1 => input_p1_times_b1_mul_componentxUMxa3_and_b4
                           , B0 => n2639, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b2, Y => 
                           n2640);
   U3162 : INVX1 port map( A => n2870, Y => n1142);
   U3163 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b2
                           , A1 => input_p2_times_b2_mul_componentxUMxa3_and_b3
                           , B0 => n2869, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b1, Y => 
                           n2870);
   U3164 : INVX1 port map( A => n3338, Y => n665);
   U3165 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b2, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b3, B0 =>
                           n3337, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b1, Y => 
                           n3338);
   U3166 : INVX1 port map( A => n2408, Y => n787);
   U3167 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b7, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b8, B0 
                           => n2407, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b6, Y => 
                           n2408);
   U3168 : INVX1 port map( A => n2406, Y => n818);
   U3169 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b3, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b4, B0 
                           => n2405, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b2, Y => 
                           n2406);
   U3170 : INVX1 port map( A => n2650, Y => n963);
   U3171 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b5
                           , A1 => input_p1_times_b1_mul_componentxUMxa3_and_b6
                           , B0 => n2649, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b4, Y => 
                           n2650);
   U3172 : INVX1 port map( A => n2968, Y => n1104);
   U3173 : AOI22X1 port map( A0 => n1105, A1 => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b0, B0 => 
                           n2967, B1 => n1128, Y => n2968);
   U3174 : INVX1 port map( A => n2884, Y => n1122);
   U3175 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b5
                           , A1 => input_p2_times_b2_mul_componentxUMxa3_and_b6
                           , B0 => n2883, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b4, Y => 
                           n2884);
   U3176 : INVX1 port map( A => n3436, Y => n627);
   U3177 : AOI22X1 port map( A0 => n628, A1 => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b0, B0 =>
                           n3435, B1 => n651, Y => n3436);
   U3178 : INVX1 port map( A => n3352, Y => n645);
   U3179 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b5, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b6, B0 =>
                           n3351, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b4, Y => 
                           n3352);
   U3180 : INVX1 port map( A => n2416, Y => n804);
   U3181 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b5, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b6, B0 
                           => n2415, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b4, Y => 
                           n2416);
   U3182 : INVX1 port map( A => n2890, Y => n1112);
   U3183 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b6
                           , A1 => input_p2_times_b2_mul_componentxUMxa3_and_b7
                           , B0 => n2889, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b5, Y => 
                           n2890);
   U3184 : INVX1 port map( A => n3358, Y => n635);
   U3185 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b6, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b7, B0 =>
                           n3357, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b5, Y => 
                           n3358);
   U3186 : INVX1 port map( A => n2908, Y => n1140);
   U3187 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b2, A1 =>
                           input_p2_times_b2_mul_componentxUMxa9_and_b3, B0 => 
                           n2907, B1 => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b1, Y => 
                           n2908);
   U3188 : INVX1 port map( A => n3376, Y => n663);
   U3189 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b2, A1 
                           => output_p2_times_a2_mul_componentxUMxa9_and_b3, B0
                           => n3375, B1 => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b1, Y =>
                           n3376);
   U3190 : INVX1 port map( A => n2916, Y => n1134);
   U3191 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b3, A1 =>
                           input_p2_times_b2_mul_componentxUMxa9_and_b4, B0 => 
                           n2915, B1 => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b2, Y => 
                           n2916);
   U3192 : INVX1 port map( A => n3384, Y => n657);
   U3193 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b3, A1 
                           => output_p2_times_a2_mul_componentxUMxa9_and_b4, B0
                           => n3383, B1 => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b2, Y =>
                           n3384);
   U3194 : INVX1 port map( A => n2746, Y => n911);
   U3195 : AOI22X1 port map( A0 => n912, A1 => 
                           input_p1_times_b1_mul_componentxUMxa12_and_b0, B0 =>
                           n2745, B1 => n944, Y => n2746);
   U3196 : INVX1 port map( A => n2980, Y => n1070);
   U3197 : AOI22X1 port map( A0 => n1071, A1 => 
                           input_p2_times_b2_mul_componentxUMxa12_and_b0, B0 =>
                           n2979, B1 => n1103, Y => n2980);
   U3198 : INVX1 port map( A => n3448, Y => n593);
   U3199 : AOI22X1 port map( A0 => n594, A1 => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b0, B0 
                           => n3447, B1 => n626, Y => n3448);
   U3200 : INVX1 port map( A => n2512, Y => n752);
   U3201 : AOI22X1 port map( A0 => n753, A1 => 
                           input_times_b0_mul_componentxUMxa12_and_b0, B0 => 
                           n2511, B1 => n785, Y => n2512);
   U3202 : INVX1 port map( A => n2626, Y => n985);
   U3203 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b2
                           , A1 => input_p1_times_b1_mul_componentxUMxa0_and_b3
                           , B0 => n2625, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b1, Y => 
                           n2626);
   U3204 : INVX1 port map( A => n2392, Y => n826);
   U3205 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b2, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b3, B0 
                           => n2391, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b1, Y => 
                           n2392);
   U3206 : INVX1 port map( A => n2634, Y => n964);
   U3207 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b5
                           , A1 => input_p1_times_b1_mul_componentxUMxa0_and_b6
                           , B0 => n2633, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b4, Y => 
                           n2634);
   U3208 : INVX1 port map( A => n2638, Y => n956);
   U3209 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b6
                           , A1 => input_p1_times_b1_mul_componentxUMxa0_and_b7
                           , B0 => n2637, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b5, Y => 
                           n2638);
   U3210 : INVX1 port map( A => n2868, Y => n1123);
   U3211 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b5
                           , A1 => input_p2_times_b2_mul_componentxUMxa0_and_b6
                           , B0 => n2867, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b4, Y => 
                           n2868);
   U3212 : INVX1 port map( A => n3336, Y => n646);
   U3213 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b5, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b6, B0 =>
                           n3335, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b4, Y => 
                           n3336);
   U3214 : INVX1 port map( A => n2400, Y => n805);
   U3215 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b5, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b6, B0 
                           => n2399, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b4, Y => 
                           n2400);
   U3216 : INVX1 port map( A => n2404, Y => n797);
   U3217 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b6, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b7, B0 
                           => n2403, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b5, Y => 
                           n2404);
   U3218 : INVX1 port map( A => n2880, Y => n1148);
   U3219 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b1
                           , A1 => input_p2_times_b2_mul_componentxUMxa6_and_b2
                           , B0 => n2879, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b0, Y => 
                           n2880);
   U3220 : INVX1 port map( A => n3348, Y => n671);
   U3221 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b1, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b2, B0 =>
                           n3347, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b0, Y => 
                           n3348);
   U3222 : INVX1 port map( A => n2692, Y => n991);
   U3223 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa13_and_b1, A1 =>
                           input_p1_times_b1_mul_componentxUMxa12_and_b2, B0 =>
                           n2691, B1 => 
                           input_p1_times_b1_mul_componentxUMxa14_and_b0, Y => 
                           n2692);
   U3224 : INVX1 port map( A => n2926, Y => n1150);
   U3225 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa13_and_b1, A1 =>
                           input_p2_times_b2_mul_componentxUMxa12_and_b2, B0 =>
                           n2925, B1 => 
                           input_p2_times_b2_mul_componentxUMxa14_and_b0, Y => 
                           n2926);
   U3226 : INVX1 port map( A => n3394, Y => n673);
   U3227 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b1, A1 
                           => output_p2_times_a2_mul_componentxUMxa12_and_b2, 
                           B0 => n3393, B1 => 
                           output_p2_times_a2_mul_componentxUMxa14_and_b0, Y =>
                           n3394);
   U3228 : INVX1 port map( A => n2458, Y => n832);
   U3229 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa13_and_b1, 
                           A1 => input_times_b0_mul_componentxUMxa12_and_b2, B0
                           => n2457, B1 => 
                           input_times_b0_mul_componentxUMxa14_and_b0, Y => 
                           n2458);
   U3230 : INVX1 port map( A => n2632, Y => n990);
   U3231 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b1
                           , A1 => input_p1_times_b1_mul_componentxUMxa3_and_b2
                           , B0 => n2631, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b0, Y => 
                           n2632);
   U3232 : INVX1 port map( A => n2866, Y => n1149);
   U3233 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b1
                           , A1 => input_p2_times_b2_mul_componentxUMxa3_and_b2
                           , B0 => n2865, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b0, Y => 
                           n2866);
   U3234 : INVX1 port map( A => n3334, Y => n672);
   U3235 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b1, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b2, B0 =>
                           n3333, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b0, Y => 
                           n3334);
   U3236 : INVX1 port map( A => n2398, Y => n831);
   U3237 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b1, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b2, B0 
                           => n2397, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b0, Y => 
                           n2398);
   U3238 : INVX1 port map( A => n2644, Y => n969);
   U3239 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b4
                           , A1 => input_p1_times_b1_mul_componentxUMxa3_and_b5
                           , B0 => n2643, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b3, Y => 
                           n2644);
   U3240 : INVX1 port map( A => n2878, Y => n1128);
   U3241 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b4
                           , A1 => input_p2_times_b2_mul_componentxUMxa3_and_b5
                           , B0 => n2877, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b3, Y => 
                           n2878);
   U3242 : INVX1 port map( A => n3346, Y => n651);
   U3243 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b4, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b5, B0 =>
                           n3345, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b3, Y => 
                           n3346);
   U3244 : INVX1 port map( A => n2410, Y => n810);
   U3245 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b4, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b5, B0 
                           => n2409, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b3, Y => 
                           n2410);
   U3246 : INVX1 port map( A => n2652, Y => n982);
   U3247 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b2
                           , A1 => input_p1_times_b1_mul_componentxUMxa6_and_b3
                           , B0 => n2651, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b1, Y => 
                           n2652);
   U3248 : INVX1 port map( A => n2886, Y => n1141);
   U3249 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b2
                           , A1 => input_p2_times_b2_mul_componentxUMxa6_and_b3
                           , B0 => n2885, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b1, Y => 
                           n2886);
   U3250 : INVX1 port map( A => n3354, Y => n664);
   U3251 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b2, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b3, B0 =>
                           n3353, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b1, Y => 
                           n3354);
   U3252 : INVX1 port map( A => n2418, Y => n823);
   U3253 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b2, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b3, B0 
                           => n2417, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b1, Y => 
                           n2418);
   U3254 : INVX1 port map( A => n2658, Y => n976);
   U3255 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b3
                           , A1 => input_p1_times_b1_mul_componentxUMxa6_and_b4
                           , B0 => n2657, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b2, Y => 
                           n2658);
   U3256 : INVX1 port map( A => n2892, Y => n1135);
   U3257 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b3
                           , A1 => input_p2_times_b2_mul_componentxUMxa6_and_b4
                           , B0 => n2891, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b2, Y => 
                           n2892);
   U3258 : INVX1 port map( A => n3360, Y => n658);
   U3259 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b3, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b4, B0 =>
                           n3359, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b2, Y => 
                           n3360);
   U3260 : INVX1 port map( A => n2424, Y => n817);
   U3261 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b3, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b4, B0 
                           => n2423, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b2, Y => 
                           n2424);
   U3262 : INVX1 port map( A => n2700, Y => n961);
   U3263 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b5, A1 =>
                           input_p1_times_b1_mul_componentxUMxa9_and_b6, B0 => 
                           n2699, B1 => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b4, Y => 
                           n2700);
   U3264 : INVX1 port map( A => n2466, Y => n802);
   U3265 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa10_and_b5, 
                           A1 => input_times_b0_mul_componentxUMxa9_and_b6, B0 
                           => n2465, B1 => 
                           input_times_b0_mul_componentxUMxa11_and_b4, Y => 
                           n2466);
   U3266 : INVX1 port map( A => n2912, Y => n1082);
   U3267 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b9
                           , A1 => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b10, B0 =>
                           n2911, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b8, Y => 
                           n2912);
   U3268 : INVX1 port map( A => n3380, Y => n605);
   U3269 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b9, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b10, B0 
                           => n3379, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b8, Y => 
                           n3380);
   U3270 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa13_and_b3, A1 =>
                           input_p1_times_b1_mul_componentxUMxa12_and_b4, B0 =>
                           n2711, B1 => 
                           input_p1_times_b1_mul_componentxUMxa14_and_b2, Y => 
                           n2712);
   U3271 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa13_and_b3, A1 =>
                           input_p2_times_b2_mul_componentxUMxa12_and_b4, B0 =>
                           n2945, B1 => 
                           input_p2_times_b2_mul_componentxUMxa14_and_b2, Y => 
                           n2946);
   U3272 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b3, A1 
                           => output_p2_times_a2_mul_componentxUMxa12_and_b4, 
                           B0 => n3413, B1 => 
                           output_p2_times_a2_mul_componentxUMxa14_and_b2, Y =>
                           n3414);
   U3273 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa13_and_b3, 
                           A1 => input_times_b0_mul_componentxUMxa12_and_b4, B0
                           => n2477, B1 => 
                           input_times_b0_mul_componentxUMxa14_and_b2, Y => 
                           n2478);
   U3274 : INVX1 port map( A => n2882, Y => n1094);
   U3275 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b8
                           , A1 => input_p2_times_b2_mul_componentxUMxa0_and_b9
                           , B0 => n2881, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b7, Y => 
                           n2882);
   U3276 : INVX1 port map( A => n2904, Y => n1091);
   U3277 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b8
                           , A1 => input_p2_times_b2_mul_componentxUMxa3_and_b9
                           , B0 => n2903, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b7, Y => 
                           n2904);
   U3278 : INVX1 port map( A => n3350, Y => n617);
   U3279 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b8, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b9, B0 =>
                           n3349, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b7, Y => 
                           n3350);
   U3280 : INVX1 port map( A => n3372, Y => n614);
   U3281 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b8, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b9, B0 =>
                           n3371, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b7, Y => 
                           n3372);
   U3282 : INVX1 port map( A => n2922, Y => n1102);
   U3283 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b7
                           , A1 => input_p2_times_b2_mul_componentxUMxa6_and_b8
                           , B0 => n2921, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b6, Y => 
                           n2922);
   U3284 : INVX1 port map( A => n3390, Y => n625);
   U3285 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b7, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b8, B0 =>
                           n3389, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b6, Y => 
                           n3390);
   U3286 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b11,
                           B => n2675, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831568_127845824_127847728);
   U3287 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b11,
                           B => n2909, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831568_127845824_127847728);
   U3288 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b11
                           , B => n3377, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831568_127845824_127847728);
   U3289 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b11, B 
                           => n2441, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831568_127845824_127847728);
   U3290 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b7, 
                           B => n2647, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831120_127845376_127847280);
   U3291 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b7, 
                           B => n2881, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831120_127845376_127847280);
   U3292 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b7,
                           B => n3349, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831120_127845376_127847280);
   U3293 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b7, B 
                           => n2413, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831120_127845376_127847280);
   U3294 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b9, 
                           B => n2659, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831344_127845600_127847504);
   U3295 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b9, 
                           B => n2893, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831344_127845600_127847504);
   U3296 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b9,
                           B => n3361, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831344_127845600_127847504);
   U3297 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b9, B 
                           => n2425, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831344_127845600_127847504);
   U3298 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b6, 
                           B => n2921, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732704_127722384_127724288);
   U3299 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b6,
                           B => n3389, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732704_127722384_127724288);
   U3300 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b10,
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b9, Y
                           => n2653);
   U3301 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b10,
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b9, Y
                           => n2887);
   U3302 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b10
                           , B => output_p2_times_a2_mul_componentxUMxa1_and_b9
                           , Y => n3355);
   U3303 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b10, B 
                           => input_times_b0_mul_componentxUMxa1_and_b9, Y => 
                           n2419);
   U3304 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b10,
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b9, Y
                           => n2677);
   U3305 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b10,
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b9, Y
                           => n2911);
   U3306 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b10
                           , B => output_p2_times_a2_mul_componentxUMxa4_and_b9
                           , Y => n3379);
   U3307 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b10, B 
                           => input_times_b0_mul_componentxUMxa4_and_b9, Y => 
                           n2443);
   U3308 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b11,
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b10, 
                           Y => n2685);
   U3309 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b11,
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b10, 
                           Y => n2919);
   U3310 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b11
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b10, Y =>
                           n3387);
   U3311 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b11, B 
                           => input_times_b0_mul_componentxUMxa4_and_b10, Y => 
                           n2451);
   U3312 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b11,
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b10, 
                           Y => n2659);
   U3313 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b11,
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b10, 
                           Y => n2893);
   U3314 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b11
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b10, Y =>
                           n3361);
   U3315 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b11, B 
                           => input_times_b0_mul_componentxUMxa1_and_b10, Y => 
                           n2425);
   U3316 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa12_and_b4,
                           B => input_p1_times_b1_mul_componentxUMxa13_and_b3, 
                           Y => n2711);
   U3317 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa12_and_b4, B 
                           => input_times_b0_mul_componentxUMxa13_and_b3, Y => 
                           n2477);
   U3318 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b12,
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b11, 
                           Y => n2667);
   U3319 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b12,
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b11, 
                           Y => n2901);
   U3320 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b12
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b11, Y =>
                           n3369);
   U3321 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b12, B 
                           => input_times_b0_mul_componentxUMxa1_and_b11, Y => 
                           n2433);
   U3322 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa12_and_b4,
                           B => input_p2_times_b2_mul_componentxUMxa13_and_b3, 
                           Y => n2945);
   U3323 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa12_and_b4
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b3, Y =>
                           n3413);
   U3324 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b13,
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b12, 
                           Y => n2675);
   U3325 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b13,
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b12, 
                           Y => n2909);
   U3326 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b13
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b12, Y =>
                           n3377);
   U3327 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b13, B 
                           => input_times_b0_mul_componentxUMxa1_and_b12, Y => 
                           n2441);
   U3328 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b2, 
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b1, Y
                           => n2623);
   U3329 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b2, 
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b1, Y
                           => n2857);
   U3330 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b2,
                           B => output_p2_times_a2_mul_componentxUMxa1_and_b1, 
                           Y => n3325);
   U3331 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b2, B 
                           => input_times_b0_mul_componentxUMxa1_and_b1, Y => 
                           input_times_b0_mul_componentxUMxFA_127826296_127826240xn2);
   U3332 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b9, 
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b8, Y
                           => n2647);
   U3333 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b9, 
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b8, Y
                           => n2881);
   U3334 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b9,
                           B => output_p2_times_a2_mul_componentxUMxa1_and_b8, 
                           Y => n3349);
   U3335 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b9, B 
                           => input_times_b0_mul_componentxUMxa1_and_b8, Y => 
                           n2413);
   U3336 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b0, 
                           B => n992, Y => n2719);
   U3337 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b0, 
                           B => n1151, Y => n2953);
   U3338 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b0,
                           B => n674, Y => n3421);
   U3339 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b0, B 
                           => n833, Y => n2485);
   U3340 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b9, 
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b8, Y
                           => n2669);
   U3341 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b9, 
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b8, Y
                           => n2903);
   U3342 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b9,
                           B => output_p2_times_a2_mul_componentxUMxa4_and_b8, 
                           Y => n3371);
   U3343 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b9, B 
                           => input_times_b0_mul_componentxUMxa4_and_b8, Y => 
                           n2435);
   U3344 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b8, 
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b7, Y
                           => n2661);
   U3345 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b8, 
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b7, Y
                           => n2895);
   U3346 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b8,
                           B => output_p2_times_a2_mul_componentxUMxa4_and_b7, 
                           Y => n3363);
   U3347 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b8, B 
                           => input_times_b0_mul_componentxUMxa4_and_b7, Y => 
                           n2427);
   U3348 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b7, 
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b6, Y
                           => n2679);
   U3349 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b7, 
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b6, Y
                           => n2913);
   U3350 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b7,
                           B => output_p2_times_a2_mul_componentxUMxa7_and_b6, 
                           Y => n3381);
   U3351 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b7, B 
                           => input_times_b0_mul_componentxUMxa7_and_b6, Y => 
                           n2445);
   U3352 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b8, 
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b7, Y
                           => n2921);
   U3353 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b8,
                           B => output_p2_times_a2_mul_componentxUMxa7_and_b7, 
                           Y => n3389);
   U3354 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa9_and_b6, 
                           B => input_p1_times_b1_mul_componentxUMxa10_and_b5, 
                           Y => n2699);
   U3355 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b9, 
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b8, Y
                           => n2697);
   U3356 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa9_and_b6, 
                           B => input_p2_times_b2_mul_componentxUMxa10_and_b5, 
                           Y => n2933);
   U3357 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa9_and_b6,
                           B => output_p2_times_a2_mul_componentxUMxa10_and_b5,
                           Y => n3401);
   U3358 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa9_and_b6, B 
                           => input_times_b0_mul_componentxUMxa10_and_b5, Y => 
                           n2465);
   U3359 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b9, B 
                           => input_times_b0_mul_componentxUMxa7_and_b8, Y => 
                           n2463);
   U3360 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa9_and_b7, 
                           B => input_p1_times_b1_mul_componentxUMxa10_and_b6, 
                           Y => n2709);
   U3361 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa9_and_b7, 
                           B => input_p2_times_b2_mul_componentxUMxa10_and_b6, 
                           Y => n2943);
   U3362 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa9_and_b7,
                           B => output_p2_times_a2_mul_componentxUMxa10_and_b6,
                           Y => n3411);
   U3363 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa9_and_b7, B 
                           => input_times_b0_mul_componentxUMxa10_and_b6, Y => 
                           n2475);
   U3364 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b0, 
                           B => n2631, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672672_127674576_127729792);
   U3365 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b0, 
                           B => n2865, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672672_127674576_127729792);
   U3366 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b0,
                           B => n3333, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672672_127674576_127729792);
   U3367 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b0, B 
                           => n2397, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672672_127674576_127729792);
   U3368 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b5, 
                           B => n2679, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732592_127722272_127724176);
   U3369 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b5, 
                           B => n2913, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732592_127722272_127724176);
   U3370 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b5,
                           B => n3381, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732592_127722272_127724176);
   U3371 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b5, B 
                           => n2445, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732592_127722272_127724176);
   U3372 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b8, 
                           B => n2653, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831232_127845488_127847392);
   U3373 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b8, 
                           B => n2887, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831232_127845488_127847392);
   U3374 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b8,
                           B => n3355, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831232_127845488_127847392);
   U3375 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b8, B 
                           => n2419, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831232_127845488_127847392);
   U3376 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b7, 
                           B => n2669, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673456_127675360_127730576);
   U3377 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b7, 
                           B => n2903, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673456_127675360_127730576);
   U3378 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b7,
                           B => n3371, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673456_127675360_127730576);
   U3379 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b7, B 
                           => n2435, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673456_127675360_127730576);
   U3380 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b9, 
                           B => n2685, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673680_127675584_127730800);
   U3381 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b9, 
                           B => n2919, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673680_127675584_127730800);
   U3382 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b9,
                           B => n3387, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673680_127675584_127730800);
   U3383 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b9, B 
                           => n2451, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673680_127675584_127730800);
   U3384 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b10,
                           B => n2667, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831456_127845712_127847616);
   U3385 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b10,
                           B => n2901, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831456_127845712_127847616);
   U3386 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b10
                           , B => n3369, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831456_127845712_127847616);
   U3387 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b10, B 
                           => n2433, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831456_127845712_127847616);
   U3388 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa11_and_b5,
                           B => n2709, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636368_127638272_127713968);
   U3389 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa11_and_b5, B 
                           => n2475, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636368_127638272_127713968);
   U3390 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa11_and_b5,
                           B => n2943, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636368_127638272_127713968);
   U3391 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa11_and_b5
                           , B => n3411, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636368_127638272_127713968);
   U3392 : OAI2BB2X1 port map( B0 => n133, B1 => n1260, A0N => 
                           output_previous_2_17_port, A1N => n319, Y => n4672);
   U3393 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b1, 
                           B => n2625, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830448_127844704_127846608);
   U3394 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b1, 
                           B => n2859, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830448_127844704_127846608);
   U3395 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b1,
                           B => n3327, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830448_127844704_127846608);
   U3396 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b1, B 
                           => n2391, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830448_127844704_127846608);
   U3397 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b4, 
                           B => n2883, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673120_127675024_127730240);
   U3398 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b4,
                           B => n3351, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673120_127675024_127730240);
   U3399 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b6, 
                           B => n2661, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673344_127675248_127730464);
   U3400 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b6, 
                           B => n2895, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673344_127675248_127730464);
   U3401 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b6,
                           B => n3363, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673344_127675248_127730464);
   U3402 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b6, B 
                           => n2427, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673344_127675248_127730464);
   U3403 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b7, 
                           B => n2697, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732816_127722496_127724400);
   U3404 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b7, B 
                           => n2463, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732816_127722496_127724400);
   U3405 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b8, 
                           B => n2677, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673568_127675472_127730688);
   U3406 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b8, 
                           B => n2911, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673568_127675472_127730688);
   U3407 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b8,
                           B => n3379, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673568_127675472_127730688);
   U3408 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b8, B 
                           => n2443, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673568_127675472_127730688);
   U3409 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa4_and_b0, 
                           B => input_p1_times_b1_mul_componentxUMxa3_and_b1, Y
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127672560_127674464);
   U3410 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa4_and_b0, 
                           B => input_p2_times_b2_mul_componentxUMxa3_and_b1, Y
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127672560_127674464);
   U3411 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa4_and_b0,
                           B => output_p2_times_a2_mul_componentxUMxa3_and_b1, 
                           Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127672560_127674464);
   U3412 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa4_and_b0, B 
                           => input_times_b0_mul_componentxUMxa3_and_b1, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127672560_127674464);
   U3413 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa11_and_b4,
                           B => n2699, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636256_127638160_127713856);
   U3414 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa11_and_b4, B 
                           => n2465, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636256_127638160_127713856);
   U3415 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa11_and_b4,
                           B => n2933, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636256_127638160_127713856);
   U3416 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa11_and_b4
                           , B => n3401, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636256_127638160_127713856);
   U3417 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa14_and_b2,
                           B => n2711, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715872_127848912_127850816);
   U3418 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa14_and_b2, B 
                           => n2477, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715872_127848912_127850816);
   U3419 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa14_and_b2,
                           B => n2945, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715872_127848912_127850816);
   U3420 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa14_and_b2
                           , B => n3413, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715872_127848912_127850816);
   U3421 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b3, 
                           B => n2663, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732368_127722048_127723952);
   U3422 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b3, 
                           B => n2897, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732368_127722048_127723952);
   U3423 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b3,
                           B => n3365, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732368_127722048_127723952);
   U3424 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b3, B 
                           => n2429, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732368_127722048_127723952);
   U3425 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa14_and_b1,
                           B => n2701, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715760_127848800_127850704);
   U3426 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa14_and_b1, B 
                           => n2467, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715760_127848800_127850704);
   U3427 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa14_and_b1,
                           B => n2935, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715760_127848800_127850704);
   U3428 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa14_and_b1
                           , B => n3403, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715760_127848800_127850704);
   U3429 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b0, 
                           B => n2623, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830336_127844592_127846496);
   U3430 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b0, 
                           B => n2857, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830336_127844592_127846496);
   U3431 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b0,
                           B => n3325, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830336_127844592_127846496);
   U3432 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b0, B 
                           => 
                           input_times_b0_mul_componentxUMxFA_127826296_127826240xn2, Y 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830336_127844592_127846496);
   U3433 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa16_and_b0,
                           B => input_p1_times_b1_mul_componentxUMxa15_and_b1, 
                           Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127627504_127629408);
   U3434 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa16_and_b0, B 
                           => input_times_b0_mul_componentxUMxa15_and_b1, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127627504_127629408);
   U3435 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa16_and_b0,
                           B => input_p2_times_b2_mul_componentxUMxa15_and_b1, 
                           Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127627504_127629408);
   U3436 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa16_and_b0
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa15_and_b1, Y =>
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127627504_127629408);
   U3437 : XOR2X1 port map( A => n2710, B => n2712, Y => n2776);
   U3438 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b6, A1 =>
                           input_p1_times_b1_mul_componentxUMxa9_and_b7, B0 => 
                           n2709, B1 => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b5, Y => 
                           n2710);
   U3439 : XOR2X1 port map( A => n2944, B => n2946, Y => n3010);
   U3440 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b6, A1 =>
                           input_p2_times_b2_mul_componentxUMxa9_and_b7, B0 => 
                           n2943, B1 => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b5, Y => 
                           n2944);
   U3441 : XOR2X1 port map( A => n3412, B => n3414, Y => n3478);
   U3442 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b6, A1 
                           => output_p2_times_a2_mul_componentxUMxa9_and_b7, B0
                           => n3411, B1 => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b5, Y =>
                           n3412);
   U3443 : XOR2X1 port map( A => n2476, B => n2478, Y => n2542);
   U3444 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa10_and_b6, 
                           A1 => input_times_b0_mul_componentxUMxa9_and_b7, B0 
                           => n2475, B1 => 
                           input_times_b0_mul_componentxUMxa11_and_b5, Y => 
                           n2476);
   U3445 : INVX1 port map( A => n2660, Y => n912);
   U3446 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b10, A1 =>
                           input_p1_times_b1_mul_componentxUMxa0_and_b11, B0 =>
                           n2659, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b9, Y => 
                           n2660);
   U3447 : INVX1 port map( A => n2894, Y => n1071);
   U3448 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b10, A1 =>
                           input_p2_times_b2_mul_componentxUMxa0_and_b11, B0 =>
                           n2893, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b9, Y => 
                           n2894);
   U3449 : INVX1 port map( A => n3362, Y => n594);
   U3450 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b10, A1 
                           => output_p2_times_a2_mul_componentxUMxa0_and_b11, 
                           B0 => n3361, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b9, Y => 
                           n3362);
   U3451 : INVX1 port map( A => n2426, Y => n753);
   U3452 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b10, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b11, B0
                           => n2425, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b9, Y => 
                           n2426);
   U3453 : INVX1 port map( A => n2678, Y => n923);
   U3454 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b9
                           , A1 => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b10, B0 =>
                           n2677, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b8, Y => 
                           n2678);
   U3455 : INVX1 port map( A => n2444, Y => n764);
   U3456 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b9, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b10, B0
                           => n2443, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b8, Y => 
                           n2444);
   U3457 : INVX1 port map( A => n2876, Y => n1105);
   U3458 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b7
                           , A1 => input_p2_times_b2_mul_componentxUMxa0_and_b8
                           , B0 => n2875, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b6, Y => 
                           n2876);
   U3459 : INVX1 port map( A => n3344, Y => n628);
   U3460 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b7, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b8, B0 =>
                           n3343, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b6, Y => 
                           n3344);
   U3461 : INVX1 port map( A => n2624, Y => n992);
   U3462 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b1
                           , A1 => input_p1_times_b1_mul_componentxUMxa0_and_b2
                           , B0 => n2623, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b0, Y => 
                           n2624);
   U3463 : INVX1 port map( A => n2858, Y => n1151);
   U3464 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b1
                           , A1 => input_p2_times_b2_mul_componentxUMxa0_and_b2
                           , B0 => n2857, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b0, Y => 
                           n2858);
   U3465 : INVX1 port map( A => n3326, Y => n674);
   U3466 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b1, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b2, B0 =>
                           n3325, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b0, Y => 
                           n3326);
   U3467 : INVX1 port map( A => 
                           input_times_b0_mul_componentxUMxFA_127826296_127826240xn3, Y 
                           => n833);
   U3468 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b1, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b2, B0 
                           => 
                           input_times_b0_mul_componentxUMxFA_127826296_127826240xn2, 
                           B1 => input_times_b0_mul_componentxUMxa2_and_b0, Y 
                           => 
                           input_times_b0_mul_componentxUMxFA_127826296_127826240xn3);
   U3469 : INVX1 port map( A => n2670, Y => n932);
   U3470 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b8
                           , A1 => input_p1_times_b1_mul_componentxUMxa3_and_b9
                           , B0 => n2669, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b7, Y => 
                           n2670);
   U3471 : INVX1 port map( A => n2436, Y => n773);
   U3472 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b8, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b9, B0 
                           => n2435, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b7, Y => 
                           n2436);
   U3473 : INVX1 port map( A => n2654, Y => n927);
   U3474 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b9
                           , A1 => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b10, B0 =>
                           n2653, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b8, Y => 
                           n2654);
   U3475 : INVX1 port map( A => n2888, Y => n1086);
   U3476 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa1_and_b9
                           , A1 => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b10, B0 =>
                           n2887, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b8, Y => 
                           n2888);
   U3477 : INVX1 port map( A => n3356, Y => n609);
   U3478 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b9, A1 =>
                           output_p2_times_a2_mul_componentxUMxa0_and_b10, B0 
                           => n3355, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b8, Y => 
                           n3356);
   U3479 : INVX1 port map( A => n2420, Y => n768);
   U3480 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b9, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b10, B0
                           => n2419, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b8, Y => 
                           n2420);
   U3481 : INVX1 port map( A => n2668, Y => n904);
   U3482 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b11, A1 =>
                           input_p1_times_b1_mul_componentxUMxa0_and_b12, B0 =>
                           n2667, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b10, Y => 
                           n2668);
   U3483 : INVX1 port map( A => n2902, Y => n1063);
   U3484 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b11, A1 =>
                           input_p2_times_b2_mul_componentxUMxa0_and_b12, B0 =>
                           n2901, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b10, Y => 
                           n2902);
   U3485 : INVX1 port map( A => n3370, Y => n586);
   U3486 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b11, A1 
                           => output_p2_times_a2_mul_componentxUMxa0_and_b12, 
                           B0 => n3369, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b10, Y =>
                           n3370);
   U3487 : INVX1 port map( A => n2434, Y => n745);
   U3488 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b11, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b12, B0
                           => n2433, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b10, Y => 
                           n2434);
   U3489 : INVX1 port map( A => n2934, Y => n1120);
   U3490 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b5, A1 =>
                           input_p2_times_b2_mul_componentxUMxa9_and_b6, B0 => 
                           n2933, B1 => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b4, Y => 
                           n2934);
   U3491 : INVX1 port map( A => n3402, Y => n643);
   U3492 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b5, A1 
                           => output_p2_times_a2_mul_componentxUMxa9_and_b6, B0
                           => n3401, B1 => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b4, Y =>
                           n3402);
   U3493 : INVX1 port map( A => n2676, Y => n902);
   U3494 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b12, A1 =>
                           input_p1_times_b1_mul_componentxUMxa0_and_b13, B0 =>
                           n2675, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b11, Y => 
                           n2676);
   U3495 : INVX1 port map( A => n2910, Y => n1061);
   U3496 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b12, A1 =>
                           input_p2_times_b2_mul_componentxUMxa0_and_b13, B0 =>
                           n2909, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b11, Y => 
                           n2910);
   U3497 : INVX1 port map( A => n3378, Y => n584);
   U3498 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b12, A1 
                           => output_p2_times_a2_mul_componentxUMxa0_and_b13, 
                           B0 => n3377, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b11, Y =>
                           n3378);
   U3499 : INVX1 port map( A => n2442, Y => n743);
   U3500 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b12, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b13, B0
                           => n2441, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b11, Y => 
                           n2442);
   U3501 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127627616_127629520_127824000, B 
                           => n2778, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128199816_128200040_128199984);
   U3502 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636480_127638384_127714080, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715984_127849024_127850928, Y 
                           => n2778);
   U3503 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa17_and_b0,
                           B => n2718, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127627616_127629520_127824000);
   U3504 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa11_and_b6,
                           B => n2716, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127636480_127638384_127714080);
   U3505 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127627616_127629520_127824000, B 
                           => n3012, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128199816_128200040_128199984);
   U3506 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636480_127638384_127714080, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715984_127849024_127850928, Y 
                           => n3012);
   U3507 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa17_and_b0,
                           B => n2952, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127627616_127629520_127824000);
   U3508 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa11_and_b6,
                           B => n2950, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127636480_127638384_127714080);
   U3509 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127627616_127629520_127824000, B 
                           => n3480, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128199816_128200040_128199984);
   U3510 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636480_127638384_127714080, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715984_127849024_127850928, Y 
                           => n3480);
   U3511 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa17_and_b0
                           , B => n3420, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127627616_127629520_127824000);
   U3512 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa11_and_b6
                           , B => n3418, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127636480_127638384_127714080);
   U3513 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127627616_127629520_127824000, B 
                           => n2544, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128199816_128200040_128199984);
   U3514 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636480_127638384_127714080, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715984_127849024_127850928, Y 
                           => n2544);
   U3515 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa17_and_b0, B 
                           => n2484, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127627616_127629520_127824000);
   U3516 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa11_and_b6, B 
                           => n2482, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127636480_127638384_127714080);
   U3517 : INVX1 port map( A => n2648, Y => n935);
   U3518 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa1_and_b8
                           , A1 => input_p1_times_b1_mul_componentxUMxa0_and_b9
                           , B0 => n2647, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b7, Y => 
                           n2648);
   U3519 : INVX1 port map( A => n2414, Y => n776);
   U3520 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b8, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b9, B0 
                           => n2413, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b7, Y => 
                           n2414);
   U3521 : INVX1 port map( A => n2688, Y => n943);
   U3522 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b7
                           , A1 => input_p1_times_b1_mul_componentxUMxa6_and_b8
                           , B0 => n2687, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b6, Y => 
                           n2688);
   U3523 : INVX1 port map( A => n2454, Y => n784);
   U3524 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b7, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b8, B0 
                           => n2453, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b6, Y => 
                           n2454);
   U3525 : INVX1 port map( A => n2764, Y => n886);
   U3526 : AOI22X1 port map( A0 => n919, A1 => 
                           input_p1_times_b1_mul_componentxUMxa15_and_b0, B0 =>
                           n2763, B1 => n887, Y => n2764);
   U3527 : INVX1 port map( A => n2998, Y => n1045);
   U3528 : AOI22X1 port map( A0 => n1078, A1 => 
                           input_p2_times_b2_mul_componentxUMxa15_and_b0, B0 =>
                           n2997, B1 => n1046, Y => n2998);
   U3529 : INVX1 port map( A => n3466, Y => n568);
   U3530 : AOI22X1 port map( A0 => n601, A1 => 
                           output_p2_times_a2_mul_componentxUMxa15_and_b0, B0 
                           => n3465, B1 => n569, Y => n3466);
   U3531 : INVX1 port map( A => n2530, Y => n727);
   U3532 : AOI22X1 port map( A0 => n760, A1 => 
                           input_times_b0_mul_componentxUMxa15_and_b0, B0 => 
                           n2529, B1 => n728, Y => n2530);
   U3533 : INVX1 port map( A => n2662, Y => n944);
   U3534 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa4_and_b7
                           , A1 => input_p1_times_b1_mul_componentxUMxa3_and_b8
                           , B0 => n2661, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b6, Y => 
                           n2662);
   U3535 : INVX1 port map( A => n2672, Y => n962);
   U3536 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b5
                           , A1 => input_p1_times_b1_mul_componentxUMxa6_and_b6
                           , B0 => n2671, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b4, Y => 
                           n2672);
   U3537 : INVX1 port map( A => n2896, Y => n1103);
   U3538 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa4_and_b7
                           , A1 => input_p2_times_b2_mul_componentxUMxa3_and_b8
                           , B0 => n2895, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b6, Y => 
                           n2896);
   U3539 : INVX1 port map( A => n2906, Y => n1121);
   U3540 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b5
                           , A1 => input_p2_times_b2_mul_componentxUMxa6_and_b6
                           , B0 => n2905, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b4, Y => 
                           n2906);
   U3541 : INVX1 port map( A => n3364, Y => n626);
   U3542 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b7, A1 =>
                           output_p2_times_a2_mul_componentxUMxa3_and_b8, B0 =>
                           n3363, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b6, Y => 
                           n3364);
   U3543 : INVX1 port map( A => n3374, Y => n644);
   U3544 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b5, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b6, B0 =>
                           n3373, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b4, Y => 
                           n3374);
   U3545 : INVX1 port map( A => n2428, Y => n785);
   U3546 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b7, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b8, B0 
                           => n2427, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b6, Y => 
                           n2428);
   U3547 : INVX1 port map( A => n2438, Y => n803);
   U3548 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b5, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b6, B0 
                           => n2437, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b4, Y => 
                           n2438);
   U3549 : INVX1 port map( A => n2680, Y => n951);
   U3550 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b6
                           , A1 => input_p1_times_b1_mul_componentxUMxa6_and_b7
                           , B0 => n2679, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b5, Y => 
                           n2680);
   U3551 : INVX1 port map( A => n2914, Y => n1110);
   U3552 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b6
                           , A1 => input_p2_times_b2_mul_componentxUMxa6_and_b7
                           , B0 => n2913, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b5, Y => 
                           n2914);
   U3553 : INVX1 port map( A => n3382, Y => n633);
   U3554 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b6, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b7, B0 =>
                           n3381, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b5, Y => 
                           n3382);
   U3555 : INVX1 port map( A => n2446, Y => n792);
   U3556 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b6, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b7, B0 
                           => n2445, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b5, Y => 
                           n2446);
   U3557 : INVX1 port map( A => n2720, Y => n987);
   U3558 : AOI22X1 port map( A0 => n992, A1 => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b0, B0 => 
                           n2719, B1 => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127830448_127844704_127846608, Y 
                           => n2720);
   U3559 : INVX1 port map( A => n2954, Y => n1146);
   U3560 : AOI22X1 port map( A0 => n1151, A1 => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b0, B0 => 
                           n2953, B1 => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127830448_127844704_127846608, Y 
                           => n2954);
   U3561 : INVX1 port map( A => n3422, Y => n669);
   U3562 : AOI22X1 port map( A0 => n674, A1 => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b0, B0 =>
                           n3421, B1 => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127830448_127844704_127846608, Y 
                           => n3422);
   U3563 : INVX1 port map( A => n2486, Y => n828);
   U3564 : AOI22X1 port map( A0 => n833, A1 => 
                           input_times_b0_mul_componentxUMxa3_and_b0, B0 => 
                           n2485, B1 => 
                           input_times_b0_mul_componentxUMxsum_layer1_127830448_127844704_127846608, Y 
                           => n2486);
   U3565 : AND2X2 port map( A => input_p1_times_b1_mul_componentxUMxa16_and_b0,
                           B => input_p1_times_b1_mul_componentxUMxa15_and_b1, 
                           Y => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127627504_127629408);
   U3566 : AND2X2 port map( A => input_times_b0_mul_componentxUMxa16_and_b0, B 
                           => input_times_b0_mul_componentxUMxa15_and_b1, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127627504_127629408);
   U3567 : AND2X2 port map( A => input_p2_times_b2_mul_componentxUMxa16_and_b0,
                           B => input_p2_times_b2_mul_componentxUMxa15_and_b1, 
                           Y => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127627504_127629408);
   U3568 : AND2X2 port map( A => output_p2_times_a2_mul_componentxUMxa16_and_b0
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa15_and_b1, Y =>
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127627504_127629408);
   U3569 : INVX1 port map( A => n2696, Y => n879);
   U3570 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b11, A1 =>
                           input_p1_times_b1_mul_componentxUMxa3_and_b12, B0 =>
                           n2695, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b10, Y => 
                           n2696);
   U3571 : INVX1 port map( A => n2462, Y => n720);
   U3572 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b11, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b12, B0
                           => n2461, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b10, Y => 
                           n2462);
   U3573 : INVX1 port map( A => n2708, Y => n922);
   U3574 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b9
                           , A1 => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b10, B0 =>
                           n2707, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b8, Y => 
                           n2708);
   U3575 : INVX1 port map( A => n2474, Y => n763);
   U3576 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b9, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b10, B0
                           => n2473, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b8, Y => 
                           n2474);
   U3577 : INVX1 port map( A => n4449, Y => n993);
   U3578 : AOI22XL port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_2_port, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_2_port, 
                           B1 => n4442, Y => n4449);
   U3579 : XNOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_2_port, B 
                           => n3718, Y => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_2_port);
   U3580 : NOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_0_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_1_port, Y 
                           => n3718);
   U3581 : INVX1 port map( A => n4502, Y => n1152);
   U3582 : AOI22XL port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_2_port, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_2_port, 
                           B1 => n4495, Y => n4502);
   U3583 : XNOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_2_port, B 
                           => n3766, Y => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_2_port);
   U3584 : NOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_0_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_1_port, Y 
                           => n3766);
   U3585 : INVX1 port map( A => n4608, Y => n675);
   U3586 : AOI22XL port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_2_port, 
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_2_port, 
                           B1 => n4601, Y => n4608);
   U3587 : XNOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_2_port, B 
                           => n3862, Y => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_2_port);
   U3588 : NOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_0_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_1_port, Y 
                           => n3862);
   U3589 : INVX1 port map( A => input_times_b0_mul_componentxn98, Y => n834);
   U3590 : AOI22XL port map( A0 => 
                           input_times_b0_mul_componentxUMxfirst_vector_2_port,
                           A1 => n121, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_2_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn98);
   U3591 : XNOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_2_port,
                           B => n3670, Y => 
                           input_times_b0_mul_componentxunsigned_output_inverted_2_port);
   U3592 : NOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_0_port,
                           B => 
                           input_times_b0_mul_componentxUMxfirst_vector_1_port,
                           Y => n3670);
   U3593 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b10,
                           B => n2695, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673792_127675696_127730912);
   U3594 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b10,
                           B => n2929, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673792_127675696_127730912);
   U3595 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b10
                           , B => n3397, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673792_127675696_127730912);
   U3596 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b10, B 
                           => n2461, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673792_127675696_127730912);
   U3597 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b8, 
                           B => n2707, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127732928_127722608_127724512);
   U3598 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b8, 
                           B => n2941, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732928_127722608_127724512);
   U3599 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b8,
                           B => n3409, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732928_127722608_127724512);
   U3600 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b8, B 
                           => n2473, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127732928_127722608_127724512);
   U3601 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b10,
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b9, Y
                           => n2707);
   U3602 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b10,
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b9, Y
                           => n2941);
   U3603 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b10
                           , B => output_p2_times_a2_mul_componentxUMxa7_and_b9
                           , Y => n3409);
   U3604 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b10, B 
                           => input_times_b0_mul_componentxUMxa7_and_b9, Y => 
                           n2473);
   U3605 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b12,
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b11, 
                           Y => n2695);
   U3606 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b12,
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b11, 
                           Y => n2929);
   U3607 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b12
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b11, Y =>
                           n3397);
   U3608 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b12, B 
                           => input_times_b0_mul_componentxUMxa4_and_b11, Y => 
                           n2461);
   U3609 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b13,
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b12, 
                           Y => n2705);
   U3610 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b13,
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b12, 
                           Y => n2939);
   U3611 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b13
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b12, Y =>
                           n3407);
   U3612 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b13, B 
                           => input_times_b0_mul_componentxUMxa4_and_b12, Y => 
                           n2471);
   U3613 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b14,
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b13, 
                           Y => n2683);
   U3614 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b14,
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b13, 
                           Y => n2917);
   U3615 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b14
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b13, Y =>
                           n3385);
   U3616 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b14, B 
                           => input_times_b0_mul_componentxUMxa1_and_b13, Y => 
                           n2449);
   U3617 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b15,
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b14, 
                           Y => n2693);
   U3618 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b15,
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b14, 
                           Y => n2927);
   U3619 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b15
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b14, Y =>
                           n3395);
   U3620 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b15, B 
                           => input_times_b0_mul_componentxUMxa1_and_b14, Y => 
                           n2459);
   U3621 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b16,
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b15, 
                           Y => n2703);
   U3622 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b16,
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b15, 
                           Y => n2937);
   U3623 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b16
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b15, Y =>
                           n3405);
   U3624 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b16, B 
                           => input_times_b0_mul_componentxUMxa1_and_b15, Y => 
                           n2469);
   U3625 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b9, 
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b8, Y
                           => n2931);
   U3626 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b9,
                           B => output_p2_times_a2_mul_componentxUMxa7_and_b8, 
                           Y => n3399);
   U3627 : OR3XL port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_1_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_2_port, C 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_0_port, Y 
                           => n3717);
   U3628 : OR3XL port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_1_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_2_port, C 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_0_port, Y 
                           => n3765);
   U3629 : OR3XL port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_1_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_2_port, C 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_0_port, Y 
                           => n3861);
   U3630 : OR3XL port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_1_port,
                           B => 
                           input_times_b0_mul_componentxUMxfirst_vector_2_port,
                           C => 
                           input_times_b0_mul_componentxUMxfirst_vector_0_port,
                           Y => n3669);
   U3631 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b11,
                           B => n2705, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127673904_127675808_127731024);
   U3632 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b11,
                           B => n2939, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127673904_127675808_127731024);
   U3633 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b11
                           , B => n3407, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127673904_127675808_127731024);
   U3634 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b11, B 
                           => n2471, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127673904_127675808_127731024);
   U3635 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b13,
                           B => n2693, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831792_127846048_127847952);
   U3636 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b13,
                           B => n2927, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831792_127846048_127847952);
   U3637 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b13
                           , B => n3395, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831792_127846048_127847952);
   U3638 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b13, B 
                           => n2459, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831792_127846048_127847952);
   U3639 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b12,
                           B => n2683, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831680_127845936_127847840);
   U3640 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b12,
                           B => n2917, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831680_127845936_127847840);
   U3641 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b12
                           , B => n3385, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831680_127845936_127847840);
   U3642 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b12, B 
                           => n2449, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831680_127845936_127847840);
   U3643 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b14,
                           B => n2703, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127831904_127846160_127848064);
   U3644 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b14, B 
                           => n2469, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127831904_127846160_127848064);
   U3645 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b7, 
                           B => n2931, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127732816_127722496_127724400);
   U3646 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b7,
                           B => n3399, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127732816_127722496_127724400);
   U3647 : AND2X2 port map( A => input_p1_times_b1_mul_componentxUMxa1_and_b0, 
                           B => input_p1_times_b1_mul_componentxUMxa0_and_b1, Y
                           => 
                           input_p1_times_b1_mul_componentxUMxcarry_layer1_127830168_127844480);
   U3648 : AND2X2 port map( A => input_p2_times_b2_mul_componentxUMxa1_and_b0, 
                           B => input_p2_times_b2_mul_componentxUMxa0_and_b1, Y
                           => 
                           input_p2_times_b2_mul_componentxUMxcarry_layer1_127830168_127844480);
   U3649 : AND2X2 port map( A => output_p2_times_a2_mul_componentxUMxa1_and_b0,
                           B => output_p2_times_a2_mul_componentxUMxa0_and_b1, 
                           Y => 
                           output_p2_times_a2_mul_componentxUMxcarry_layer1_127830168_127844480);
   U3650 : AND2X2 port map( A => input_times_b0_mul_componentxUMxa1_and_b0, B 
                           => input_times_b0_mul_componentxUMxa0_and_b1, Y => 
                           input_times_b0_mul_componentxUMxcarry_layer1_127830168_127844480);
   U3651 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127733040_127722720_127724624, B 
                           => n2777, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer2_128199368_128199480_128199648);
   U3652 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127832016_127846272_127848176, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127674016_127675920_127731136, Y 
                           => n2777);
   U3653 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa8_and_b9, 
                           B => n2715, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127733040_127722720_127724624);
   U3654 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa2_and_b15,
                           B => n2713, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127832016_127846272_127848176);
   U3655 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127733040_127722720_127724624, B 
                           => n3011, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer2_128199368_128199480_128199648);
   U3656 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127832016_127846272_127848176, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127674016_127675920_127731136, Y 
                           => n3011);
   U3657 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa8_and_b9, 
                           B => n2949, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127733040_127722720_127724624);
   U3658 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b15,
                           B => n2947, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127832016_127846272_127848176);
   U3659 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127733040_127722720_127724624, B 
                           => n3479, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer2_128199368_128199480_128199648);
   U3660 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127832016_127846272_127848176, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127674016_127675920_127731136, Y 
                           => n3479);
   U3661 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa8_and_b9,
                           B => n3417, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127733040_127722720_127724624);
   U3662 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b15
                           , B => n3415, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127832016_127846272_127848176);
   U3663 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127733040_127722720_127724624, B 
                           => n2543, Y => 
                           input_times_b0_mul_componentxUMxsum_layer2_128199368_128199480_128199648);
   U3664 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxsum_layer1_127832016_127846272_127848176, B 
                           => 
                           input_times_b0_mul_componentxUMxsum_layer1_127674016_127675920_127731136, Y 
                           => n2543);
   U3665 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa8_and_b9, B 
                           => n2481, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127733040_127722720_127724624);
   U3666 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa2_and_b15, B 
                           => n2479, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127832016_127846272_127848176);
   U3667 : INVX1 port map( A => n2930, Y => n1038);
   U3668 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b11, A1 =>
                           input_p2_times_b2_mul_componentxUMxa3_and_b12, B0 =>
                           n2929, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b10, Y => 
                           n2930);
   U3669 : INVX1 port map( A => n3398, Y => n561);
   U3670 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b11, A1 
                           => output_p2_times_a2_mul_componentxUMxa3_and_b12, 
                           B0 => n3397, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b10, Y =>
                           n3398);
   U3671 : INVX1 port map( A => n2684, Y => n919);
   U3672 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b13, A1 =>
                           input_p1_times_b1_mul_componentxUMxa0_and_b14, B0 =>
                           n2683, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b12, Y => 
                           n2684);
   U3673 : INVX1 port map( A => n2918, Y => n1078);
   U3674 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b13, A1 =>
                           input_p2_times_b2_mul_componentxUMxa0_and_b14, B0 =>
                           n2917, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b12, Y => 
                           n2918);
   U3675 : INVX1 port map( A => n3386, Y => n601);
   U3676 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b13, A1 
                           => output_p2_times_a2_mul_componentxUMxa0_and_b14, 
                           B0 => n3385, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b12, Y =>
                           n3386);
   U3677 : INVX1 port map( A => n2450, Y => n760);
   U3678 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b13, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b14, B0
                           => n2449, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b12, Y => 
                           n2450);
   U3679 : INVX1 port map( A => n2694, Y => n920);
   U3680 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b14, A1 =>
                           input_p1_times_b1_mul_componentxUMxa0_and_b15, B0 =>
                           n2693, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b13, Y => 
                           n2694);
   U3681 : INVX1 port map( A => n2928, Y => n1079);
   U3682 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b14, A1 =>
                           input_p2_times_b2_mul_componentxUMxa0_and_b15, B0 =>
                           n2927, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b13, Y => 
                           n2928);
   U3683 : INVX1 port map( A => n3396, Y => n602);
   U3684 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b14, A1 
                           => output_p2_times_a2_mul_componentxUMxa0_and_b15, 
                           B0 => n3395, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b13, Y =>
                           n3396);
   U3685 : INVX1 port map( A => n2460, Y => n761);
   U3686 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b14, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b15, B0
                           => n2459, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b13, Y => 
                           n2460);
   U3687 : INVX1 port map( A => n2686, Y => n887);
   U3688 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b10, A1 =>
                           input_p1_times_b1_mul_componentxUMxa3_and_b11, B0 =>
                           n2685, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b9, Y => 
                           n2686);
   U3689 : INVX1 port map( A => n2920, Y => n1046);
   U3690 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b10, A1 =>
                           input_p2_times_b2_mul_componentxUMxa3_and_b11, B0 =>
                           n2919, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b9, Y => 
                           n2920);
   U3691 : INVX1 port map( A => n3388, Y => n569);
   U3692 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b10, A1 
                           => output_p2_times_a2_mul_componentxUMxa3_and_b11, 
                           B0 => n3387, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b9, Y => 
                           n3388);
   U3693 : INVX1 port map( A => n2452, Y => n728);
   U3694 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b10, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b11, B0
                           => n2451, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b9, Y => 
                           n2452);
   U3695 : INVX1 port map( A => n2698, Y => n931);
   U3696 : AOI22X1 port map( A0 => input_p1_times_b1_mul_componentxUMxa7_and_b8
                           , A1 => input_p1_times_b1_mul_componentxUMxa6_and_b9
                           , B0 => n2697, B1 => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b7, Y => 
                           n2698);
   U3697 : INVX1 port map( A => n2932, Y => n1090);
   U3698 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b8
                           , A1 => input_p2_times_b2_mul_componentxUMxa6_and_b9
                           , B0 => n2931, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b7, Y => 
                           n2932);
   U3699 : INVX1 port map( A => n3400, Y => n613);
   U3700 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b8, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b9, B0 =>
                           n3399, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b7, Y => 
                           n3400);
   U3701 : INVX1 port map( A => n2464, Y => n772);
   U3702 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa7_and_b8, 
                           A1 => input_times_b0_mul_componentxUMxa6_and_b9, B0 
                           => n2463, B1 => 
                           input_times_b0_mul_componentxUMxa8_and_b7, Y => 
                           n2464);
   U3703 : INVX1 port map( A => n2706, Y => n877);
   U3704 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b12, A1 =>
                           input_p1_times_b1_mul_componentxUMxa3_and_b13, B0 =>
                           n2705, B1 => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b11, Y => 
                           n2706);
   U3705 : INVX1 port map( A => n2940, Y => n1036);
   U3706 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b12, A1 =>
                           input_p2_times_b2_mul_componentxUMxa3_and_b13, B0 =>
                           n2939, B1 => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b11, Y => 
                           n2940);
   U3707 : INVX1 port map( A => n3408, Y => n559);
   U3708 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b12, A1 
                           => output_p2_times_a2_mul_componentxUMxa3_and_b13, 
                           B0 => n3407, B1 => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b11, Y =>
                           n3408);
   U3709 : INVX1 port map( A => n2472, Y => n718);
   U3710 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa4_and_b12, 
                           A1 => input_times_b0_mul_componentxUMxa3_and_b13, B0
                           => n2471, B1 => 
                           input_times_b0_mul_componentxUMxa5_and_b11, Y => 
                           n2472);
   U3711 : INVX1 port map( A => n2942, Y => n1081);
   U3712 : AOI22X1 port map( A0 => input_p2_times_b2_mul_componentxUMxa7_and_b9
                           , A1 => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b10, B0 =>
                           n2941, B1 => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b8, Y => 
                           n2942);
   U3713 : INVX1 port map( A => n3410, Y => n604);
   U3714 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b9, A1 =>
                           output_p2_times_a2_mul_componentxUMxa6_and_b10, B0 
                           => n3409, B1 => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b8, Y => 
                           n3410);
   U3715 : INVX1 port map( A => n2704, Y => n921);
   U3716 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b15, A1 =>
                           input_p1_times_b1_mul_componentxUMxa0_and_b16, B0 =>
                           n2703, B1 => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b14, Y => 
                           n2704);
   U3717 : INVX1 port map( A => n2938, Y => n1080);
   U3718 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b15, A1 =>
                           input_p2_times_b2_mul_componentxUMxa0_and_b16, B0 =>
                           n2937, B1 => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b14, Y => 
                           n2938);
   U3719 : INVX1 port map( A => n3406, Y => n603);
   U3720 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b15, A1 
                           => output_p2_times_a2_mul_componentxUMxa0_and_b16, 
                           B0 => n3405, B1 => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b14, Y =>
                           n3406);
   U3721 : INVX1 port map( A => n2470, Y => n762);
   U3722 : AOI22X1 port map( A0 => input_times_b0_mul_componentxUMxa1_and_b15, 
                           A1 => input_times_b0_mul_componentxUMxa0_and_b16, B0
                           => n2469, B1 => 
                           input_times_b0_mul_componentxUMxa2_and_b14, Y => 
                           n2470);
   U3723 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa1_and_b0, 
                           B => input_p1_times_b1_mul_componentxUMxa0_and_b1, Y
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_1_port);
   U3724 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa1_and_b0, 
                           B => input_p2_times_b2_mul_componentxUMxa0_and_b1, Y
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_1_port);
   U3725 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa1_and_b0,
                           B => output_p2_times_a2_mul_componentxUMxa0_and_b1, 
                           Y => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_1_port);
   U3726 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa1_and_b0, B 
                           => input_times_b0_mul_componentxUMxa0_and_b1, Y => 
                           input_times_b0_mul_componentxUMxfirst_vector_1_port)
                           ;
   U3727 : INVX1 port map( A => n4459, Y => n995);
   U3728 : AOI22XL port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_0_port, 
                           A1 => n125, B0 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_0_port, 
                           B1 => n4442, Y => n4459);
   U3729 : INVX1 port map( A => n4512, Y => n1154);
   U3730 : AOI22XL port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_0_port, 
                           A1 => n129, B0 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_0_port, 
                           B1 => n4495, Y => n4512);
   U3731 : INVX1 port map( A => n4618, Y => n677);
   U3732 : AOI22XL port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_0_port, 
                           A1 => n117, B0 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_0_port, 
                           B1 => n4601, Y => n4618);
   U3733 : INVX1 port map( A => input_times_b0_mul_componentxn108, Y => n836);
   U3734 : AOI22XL port map( A0 => 
                           input_times_b0_mul_componentxUMxfirst_vector_0_port,
                           A1 => n121, B0 => 
                           input_times_b0_mul_componentxUMxfirst_vector_0_port,
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn108);
   U3735 : XOR2X1 port map( A => n144, B => n334, Y => n81);
   U3736 : INVX1 port map( A => n81, Y => n4442);
   U3737 : XOR2X1 port map( A => n142, B => n325, Y => n82);
   U3738 : INVX1 port map( A => n82, Y => n4495);
   U3739 : XOR2X1 port map( A => n140, B => n352, Y => n83);
   U3740 : INVX1 port map( A => n83, Y => n4601);
   U3741 : XOR2X1 port map( A => n132, B => n343, Y => n84);
   U3742 : INVX1 port map( A => n84, Y => input_times_b0_mul_componentxn91);
   U3743 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa2_and_b14,
                           B => n2937, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127831904_127846160_127848064);
   U3744 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa2_and_b14
                           , B => n3405, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127831904_127846160_127848064);
   U3745 : INVX1 port map( A => n4450, Y => n994);
   U3746 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_1_port, 
                           A1 => n126, B0 => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_1_port, 
                           B1 => n4442, Y => n4450);
   U3747 : XOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_1_port, B 
                           => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_0_port, Y 
                           => 
                           input_p1_times_b1_mul_componentxunsigned_output_inverted_1_port);
   U3748 : INVX1 port map( A => input_times_b0_mul_componentxn99, Y => n835);
   U3749 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxUMxfirst_vector_1_port,
                           A1 => n122, B0 => 
                           input_times_b0_mul_componentxunsigned_output_inverted_1_port, 
                           B1 => input_times_b0_mul_componentxn91, Y => 
                           input_times_b0_mul_componentxn99);
   U3750 : XOR2X1 port map( A => 
                           input_times_b0_mul_componentxUMxfirst_vector_1_port,
                           B => 
                           input_times_b0_mul_componentxUMxfirst_vector_0_port,
                           Y => 
                           input_times_b0_mul_componentxunsigned_output_inverted_1_port);
   U3751 : INVX1 port map( A => n4503, Y => n1153);
   U3752 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_1_port, 
                           A1 => n130, B0 => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_1_port, 
                           B1 => n4495, Y => n4503);
   U3753 : XOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_1_port, B 
                           => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_0_port, Y 
                           => 
                           input_p2_times_b2_mul_componentxunsigned_output_inverted_1_port);
   U3754 : INVX1 port map( A => n4609, Y => n676);
   U3755 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_1_port, 
                           A1 => n118, B0 => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_1_port, 
                           B1 => n4601, Y => n4609);
   U3756 : XOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_1_port, B 
                           => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_0_port, Y 
                           => 
                           output_p2_times_a2_mul_componentxunsigned_output_inverted_1_port);
   U3757 : OAI2BB2X1 port map( B0 => n131, B1 => n319, A0N => 
                           input_previous_1_17_port, A1N => n321, Y => n4636);
   U3758 : OAI2BB2X1 port map( B0 => n143, B1 => n319, A0N => 
                           input_previous_2_17_port, A1N => n320, Y => n4654);
   U3759 : NAND3BX1 port map( AN => n845, B => input_times_b0_div_componentxn54
                           , C => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn2, Y 
                           => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn16);
   U3760 : NAND3BX1 port map( AN => n1004, B => n4232, C => n1761, Y => n1768);
   U3761 : NAND3BX1 port map( AN => n1163, B => n4288, C => n1770, Y => n1777);
   U3762 : NAND3BX1 port map( AN => n527, B => n4342, C => n1779, Y => n1786);
   U3763 : NAND3BX1 port map( AN => n686, B => n4398, C => n1788, Y => n1795);
   U3764 : NOR2BX1 port map( AN => n3892, B => parameter_B0_div(7), Y => n3891)
                           ;
   U3765 : NOR2BX1 port map( AN => n3935, B => parameter_B1_div(7), Y => n3934)
                           ;
   U3766 : NOR2BX1 port map( AN => n3978, B => parameter_B2_div(7), Y => n3977)
                           ;
   U3767 : NOR2BX1 port map( AN => n4021, B => parameter_A1_div(7), Y => n4020)
                           ;
   U3768 : NOR2BX1 port map( AN => n4064, B => parameter_A2_div(7), Y => n4063)
                           ;
   U3769 : NOR2X1 port map( A => parameter_B0_div(7), B => n3893, Y => n3892);
   U3770 : NOR2X1 port map( A => parameter_B1_div(7), B => n3936, Y => n3935);
   U3771 : NOR2X1 port map( A => parameter_B2_div(7), B => n3979, Y => n3978);
   U3772 : NOR2X1 port map( A => parameter_A1_div(7), B => n4022, Y => n4021);
   U3773 : NOR2X1 port map( A => parameter_A2_div(7), B => n4065, Y => n4064);
   U3774 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn2, B 
                           => input_times_b0_div_componentxn54, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_9_port);
   U3775 : XOR2X1 port map( A => n1761, B => n4232, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_9_port);
   U3776 : XOR2X1 port map( A => n1770, B => n4288, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_9_port);
   U3777 : XOR2X1 port map( A => n1779, B => n4342, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_9_port);
   U3778 : XOR2X1 port map( A => n1788, B => n4398, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_9_port);
   U3779 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn8, B 
                           => n849, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_3_port);
   U3780 : XOR2X1 port map( A => n1764, B => n1008, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_3_port);
   U3781 : XOR2X1 port map( A => n1773, B => n1167, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_3_port);
   U3782 : XOR2X1 port map( A => n1782, B => n531, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_3_port);
   U3783 : XOR2X1 port map( A => n1791, B => n690, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_3_port);
   U3784 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn6, B 
                           => n851, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_5_port);
   U3785 : XOR2X1 port map( A => n1763, B => n1010, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_5_port);
   U3786 : XOR2X1 port map( A => n1772, B => n1169, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_5_port);
   U3787 : XOR2X1 port map( A => n1781, B => n533, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_5_port);
   U3788 : XOR2X1 port map( A => n1790, B => n692, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_5_port);
   U3789 : OR3XL port map( A => n851, B => n852, C => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn6, Y 
                           => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn4);
   U3790 : OR3XL port map( A => n1010, B => n1011, C => n1763, Y => n1762);
   U3791 : OR3XL port map( A => n1169, B => n1170, C => n1772, Y => n1771);
   U3792 : OR3XL port map( A => n533, B => n534, C => n1781, Y => n1780);
   U3793 : OR3XL port map( A => n692, B => n693, C => n1790, Y => n1789);
   U3794 : OR2X2 port map( A => n3895, B => parameter_B0_div(7), Y => n3893);
   U3795 : OR2X2 port map( A => n3938, B => parameter_B1_div(7), Y => n3936);
   U3796 : OR2X2 port map( A => n3981, B => parameter_B2_div(7), Y => n3979);
   U3797 : OR2X2 port map( A => n4024, B => parameter_A1_div(7), Y => n4022);
   U3798 : OR2X2 port map( A => n4067, B => parameter_A2_div(7), Y => n4065);
   U3799 : XNOR2X1 port map( A => n85, B => n850, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_4_port);
   U3800 : NOR2X1 port map( A => n849, B => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn8, Y 
                           => n85);
   U3801 : XNOR2X1 port map( A => n86, B => n1009, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_4_port);
   U3802 : NOR2X1 port map( A => n1008, B => n1764, Y => n86);
   U3803 : XNOR2X1 port map( A => n87, B => n1168, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_4_port);
   U3804 : NOR2X1 port map( A => n1167, B => n1773, Y => n87);
   U3805 : XNOR2X1 port map( A => n88, B => n532, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_4_port);
   U3806 : NOR2X1 port map( A => n531, B => n1782, Y => n88);
   U3807 : XNOR2X1 port map( A => n89, B => n691, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_4_port);
   U3808 : NOR2X1 port map( A => n690, B => n1791, Y => n89);
   U3809 : XNOR2X1 port map( A => n90, B => n852, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_6_port);
   U3810 : NOR2X1 port map( A => n851, B => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn6, Y 
                           => n90);
   U3811 : XNOR2X1 port map( A => n91, B => n1011, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_6_port);
   U3812 : NOR2X1 port map( A => n1010, B => n1763, Y => n91);
   U3813 : XNOR2X1 port map( A => n92, B => n1170, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_6_port);
   U3814 : NOR2X1 port map( A => n1169, B => n1772, Y => n92);
   U3815 : XNOR2X1 port map( A => n93, B => n534, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_6_port);
   U3816 : NOR2X1 port map( A => n533, B => n1781, Y => n93);
   U3817 : XNOR2X1 port map( A => n94, B => n693, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_6_port);
   U3818 : NOR2X1 port map( A => n692, B => n1790, Y => n94);
   U3819 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn18, B 
                           => n845, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_10_port);
   U3820 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn2, B 
                           => input_times_b0_div_componentxn54, Y => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn18);
   U3821 : XOR2X1 port map( A => n1769, B => n1004, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_10_port);
   U3822 : NAND2X1 port map( A => n1761, B => n4232, Y => n1769);
   U3823 : XOR2X1 port map( A => n1778, B => n1163, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_10_port);
   U3824 : NAND2X1 port map( A => n1770, B => n4288, Y => n1778);
   U3825 : XOR2X1 port map( A => n1787, B => n527, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_10_port);
   U3826 : NAND2X1 port map( A => n1779, B => n4342, Y => n1787);
   U3827 : XOR2X1 port map( A => n1796, B => n686, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_10_port);
   U3828 : NAND2X1 port map( A => n1788, B => n4398, Y => n1796);
   U3829 : OR3XL port map( A => n849, B => n850, C => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn8, Y 
                           => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn6);
   U3830 : OR3XL port map( A => n1008, B => n1009, C => n1764, Y => n1763);
   U3831 : OR3XL port map( A => n1167, B => n1168, C => n1773, Y => n1772);
   U3832 : OR3XL port map( A => n531, B => n532, C => n1782, Y => n1781);
   U3833 : OR3XL port map( A => n690, B => n691, C => n1791, Y => n1790);
   U3834 : INVX1 port map( A => input_times_b0_div_componentxn52, Y => n853);
   U3835 : INVX1 port map( A => n4230, Y => n1012);
   U3836 : INVX1 port map( A => n4286, Y => n1171);
   U3837 : INVX1 port map( A => n4340, Y => n535);
   U3838 : INVX1 port map( A => n4396, Y => n694);
   U3839 : INVX1 port map( A => input_times_b0_div_componentxn58, Y => n840);
   U3840 : INVX1 port map( A => n4236, Y => n999);
   U3841 : INVX1 port map( A => n4292, Y => n1158);
   U3842 : INVX1 port map( A => n4346, Y => n522);
   U3843 : INVX1 port map( A => n4402, Y => n681);
   U3844 : INVX1 port map( A => input_times_b0_div_componentxn56, Y => n838);
   U3845 : INVX1 port map( A => n4234, Y => n997);
   U3846 : INVX1 port map( A => n4290, Y => n1156);
   U3847 : INVX1 port map( A => n4344, Y => n520);
   U3848 : INVX1 port map( A => n4400, Y => n679);
   U3849 : INVX1 port map( A => input_times_b0_div_componentxn53, Y => n854);
   U3850 : INVX1 port map( A => n4231, Y => n1013);
   U3851 : INVX1 port map( A => n4287, Y => n1172);
   U3852 : INVX1 port map( A => n4341, Y => n536);
   U3853 : INVX1 port map( A => n4397, Y => n695);
   U3854 : XNOR2X1 port map( A => n95, B => n843, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_16_port);
   U3855 : NOR2X1 port map( A => n842, B => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn12, Y 
                           => n95);
   U3856 : XNOR2X1 port map( A => n96, B => n1002, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_16_port);
   U3857 : NOR2X1 port map( A => n1001, B => n1766, Y => n96);
   U3858 : XNOR2X1 port map( A => n97, B => n1161, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_16_port);
   U3859 : NOR2X1 port map( A => n1160, B => n1775, Y => n97);
   U3860 : XNOR2X1 port map( A => n98, B => n525, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_16_port);
   U3861 : NOR2X1 port map( A => n524, B => n1784, Y => n98);
   U3862 : XNOR2X1 port map( A => n99, B => n684, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_16_port);
   U3863 : NOR2X1 port map( A => n683, B => n1793, Y => n99);
   U3864 : INVX1 port map( A => input_times_b0_div_componentxn57, Y => n839);
   U3865 : INVX1 port map( A => n4235, Y => n998);
   U3866 : INVX1 port map( A => n4291, Y => n1157);
   U3867 : INVX1 port map( A => n4345, Y => n521);
   U3868 : INVX1 port map( A => n4401, Y => n680);
   U3869 : INVX1 port map( A => input_times_b0_div_componentxn59, Y => n841);
   U3870 : INVX1 port map( A => n4237, Y => n1000);
   U3871 : INVX1 port map( A => n4293, Y => n1159);
   U3872 : INVX1 port map( A => n4347, Y => n523);
   U3873 : INVX1 port map( A => n4403, Y => n682);
   U3874 : INVX1 port map( A => input_times_b0_div_componentxn55, Y => n845);
   U3875 : INVX1 port map( A => n4233, Y => n1004);
   U3876 : INVX1 port map( A => n4289, Y => n1163);
   U3877 : INVX1 port map( A => n4343, Y => n527);
   U3878 : INVX1 port map( A => n4399, Y => n686);
   U3879 : INVX1 port map( A => input_times_b0_div_componentxn60, Y => n842);
   U3880 : INVX1 port map( A => n4238, Y => n1001);
   U3881 : INVX1 port map( A => n4294, Y => n1160);
   U3882 : INVX1 port map( A => n4348, Y => n524);
   U3883 : INVX1 port map( A => n4404, Y => n683);
   U3884 : INVX1 port map( A => n317, Y => n291);
   U3885 : INVX1 port map( A => n317, Y => n292);
   U3886 : INVX1 port map( A => n317, Y => n293);
   U3887 : INVX1 port map( A => n316, Y => n294);
   U3888 : INVX1 port map( A => n316, Y => n295);
   U3889 : INVX1 port map( A => n316, Y => n296);
   U3890 : INVX1 port map( A => n317, Y => n297);
   U3891 : INVX1 port map( A => reset, Y => n284);
   U3892 : INVX1 port map( A => n318, Y => n285);
   U3893 : INVX1 port map( A => n315, Y => n286);
   U3894 : INVX1 port map( A => n315, Y => n287);
   U3895 : INVX1 port map( A => n318, Y => n288);
   U3896 : INVX1 port map( A => n318, Y => n289);
   U3897 : INVX1 port map( A => n318, Y => n290);
   U3898 : INVX1 port map( A => reset, Y => n307);
   U3899 : INVX1 port map( A => reset, Y => n308);
   U3900 : INVX1 port map( A => n317, Y => n309);
   U3901 : INVX1 port map( A => n316, Y => n310);
   U3902 : INVX1 port map( A => n318, Y => n311);
   U3903 : INVX1 port map( A => n315, Y => n312);
   U3904 : INVX1 port map( A => n315, Y => n313);
   U3905 : INVX1 port map( A => n316, Y => n298);
   U3906 : INVX1 port map( A => n318, Y => n299);
   U3907 : INVX1 port map( A => n318, Y => n300);
   U3908 : INVX1 port map( A => reset, Y => n301);
   U3909 : INVX1 port map( A => n315, Y => n302);
   U3910 : INVX1 port map( A => n317, Y => n303);
   U3911 : INVX1 port map( A => n316, Y => n304);
   U3912 : INVX1 port map( A => n316, Y => n305);
   U3913 : INVX1 port map( A => n317, Y => n306);
   U3914 : INVX1 port map( A => reset, Y => n283);
   U3915 : INVX1 port map( A => n315, Y => n314);
   U3916 : AOI32X1 port map( A0 => n1320, A1 => n4135, A2 => n1340, B0 => n1311
                           , B1 => n1331, Y => n4134);
   U3917 : AOI32X1 port map( A0 => n1379, A1 => results_b0_b1_adderxn19, A2 => 
                           n1237, B0 => n1370, B1 => n1227, Y => 
                           results_b0_b1_adderxn17);
   U3918 : AOI22X1 port map( A0 => n1309, A1 => n1329, B0 => n4131, B1 => n4132
                           , Y => n4130);
   U3919 : AOI22X1 port map( A0 => n1368, A1 => n1223, B0 => 
                           results_b0_b1_adderxn14, B1 => 
                           results_b0_b1_adderxn15, Y => 
                           results_b0_b1_adderxn13);
   U3920 : AOI22X1 port map( A0 => n1307, A1 => n1327, B0 => n4127, B1 => n4128
                           , Y => n4126);
   U3921 : AOI22X1 port map( A0 => n1348, A1 => results_b0_b1_3_port, B0 => 
                           n4098, B1 => n4099, Y => n4097);
   U3922 : AOI22X1 port map( A0 => n1366, A1 => n1219, B0 => 
                           results_b0_b1_adderxn10, B1 => 
                           results_b0_b1_adderxn11, Y => results_b0_b1_adderxn9
                           );
   U3923 : AOI22X1 port map( A0 => n1305, A1 => n1325, B0 => n4123, B1 => n4124
                           , Y => n4122);
   U3924 : AOI22X1 port map( A0 => n1346, A1 => results_b0_b1_5_port, B0 => 
                           n4094, B1 => n4095, Y => n4093);
   U3925 : AOI22X1 port map( A0 => n1364, A1 => n1215, B0 => 
                           results_b0_b1_adderxn6, B1 => results_b0_b1_adderxn7
                           , Y => results_b0_b1_adderxn5);
   U3926 : AOI22X1 port map( A0 => n1344, A1 => results_b0_b1_7_port, B0 => 
                           n4090, B1 => n4091, Y => n4089);
   U3927 : AOI22X1 port map( A0 => n1362, A1 => n1211, B0 => 
                           results_b0_b1_adderxn2, B1 => results_b0_b1_adderxn3
                           , Y => results_b0_b1_adderxn34);
   U3928 : AOI22X1 port map( A0 => n1342, A1 => results_b0_b1_9_port, B0 => 
                           n4086, B1 => n4087, Y => n4117);
   U3929 : AOI22X1 port map( A0 => n1377, A1 => n1234, B0 => 
                           results_b0_b1_adderxn32, B1 => 
                           results_b0_b1_adderxn33, Y => 
                           results_b0_b1_adderxn30);
   U3930 : AOI22X1 port map( A0 => n1357, A1 => results_b0_b1_11_port, B0 => 
                           n4115, B1 => n4116, Y => n4113);
   U3931 : AOI22X1 port map( A0 => n1375, A1 => n1232, B0 => 
                           results_b0_b1_adderxn28, B1 => 
                           results_b0_b1_adderxn29, Y => 
                           results_b0_b1_adderxn26);
   U3932 : AOI22X1 port map( A0 => n1355, A1 => results_b0_b1_13_port, B0 => 
                           n4111, B1 => n4112, Y => n4109);
   U3933 : OAI2BB2X1 port map( B0 => n4101, B1 => n4100, A0N => n1349, A1N => 
                           results_b0_b1_2_port, Y => n4098);
   U3934 : OAI2BB2X1 port map( B0 => n4134, B1 => n4133, A0N => n1310, A1N => 
                           n1330, Y => n4131);
   U3935 : OAI2BB2X1 port map( B0 => results_b0_b1_adderxn17, B1 => 
                           results_b0_b1_adderxn16, A0N => n1369, A1N => n1225,
                           Y => results_b0_b1_adderxn14);
   U3936 : OAI2BB2X1 port map( B0 => n4130, B1 => n4129, A0N => n1308, A1N => 
                           n1328, Y => n4127);
   U3937 : OAI2BB2X1 port map( B0 => results_b0_b1_adderxn13, B1 => 
                           results_b0_b1_adderxn12, A0N => n1367, A1N => n1221,
                           Y => results_b0_b1_adderxn10);
   U3938 : OAI2BB2X1 port map( B0 => n4097, B1 => n4096, A0N => n1347, A1N => 
                           results_b0_b1_4_port, Y => n4094);
   U3939 : OAI2BB2X1 port map( B0 => n4126, B1 => n4125, A0N => n1306, A1N => 
                           n1326, Y => n4123);
   U3940 : OAI2BB2X1 port map( B0 => results_b0_b1_adderxn9, B1 => 
                           results_b0_b1_adderxn8, A0N => n1365, A1N => n1217, 
                           Y => results_b0_b1_adderxn6);
   U3941 : OAI2BB2X1 port map( B0 => n4093, B1 => n4092, A0N => n1345, A1N => 
                           results_b0_b1_6_port, Y => n4090);
   U3942 : OAI2BB2X1 port map( B0 => results_b0_b1_adderxn5, B1 => 
                           results_b0_b1_adderxn4, A0N => n1363, A1N => n1213, 
                           Y => results_b0_b1_adderxn2);
   U3943 : OAI2BB2X1 port map( B0 => n4089, B1 => n4088, A0N => n1343, A1N => 
                           results_b0_b1_8_port, Y => n4086);
   U3944 : OAI2BB2X1 port map( B0 => results_b0_b1_adderxn34, B1 => 
                           results_b0_b1_adderxn35, A0N => n1378, A1N => n1235,
                           Y => results_b0_b1_adderxn32);
   U3945 : OAI2BB2X1 port map( B0 => n4117, B1 => n4118, A0N => n1358, A1N => 
                           results_b0_b1_10_port, Y => n4115);
   U3946 : OAI2BB2X1 port map( B0 => results_b0_b1_adderxn30, B1 => 
                           results_b0_b1_adderxn31, A0N => n1376, A1N => n1233,
                           Y => results_b0_b1_adderxn28);
   U3947 : OAI2BB2X1 port map( B0 => n4113, B1 => n4114, A0N => n1356, A1N => 
                           results_b0_b1_12_port, Y => n4111);
   U3948 : OAI2BB2X1 port map( B0 => n4109, B1 => n4110, A0N => n1354, A1N => 
                           results_b0_b1_14_port, Y => n4107);
   U3949 : NOR2X1 port map( A => n218, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b3);
   U3950 : NOR2X1 port map( A => n217, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b4);
   U3951 : NOR2X1 port map( A => n231, B => n216, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b5);
   U3952 : XOR2X1 port map( A => results_b0_b1_3_port, B => n1348, Y => n4099);
   U3953 : XOR2X1 port map( A => results_b0_b1_5_port, B => n1346, Y => n4095);
   U3954 : XOR2X1 port map( A => results_b0_b1_7_port, B => n1344, Y => n4091);
   U3955 : XOR2X1 port map( A => results_b0_b1_9_port, B => n1342, Y => n4087);
   U3956 : XOR2X1 port map( A => results_b0_b1_11_port, B => n1357, Y => n4116)
                           ;
   U3957 : XOR2X1 port map( A => results_b0_b1_13_port, B => n1355, Y => n4112)
                           ;
   U3958 : XOR2X1 port map( A => n1331, B => n1311, Y => n4135);
   U3959 : XOR2X1 port map( A => n1227, B => n1370, Y => 
                           results_b0_b1_adderxn19);
   U3960 : XNOR2X1 port map( A => results_b0_b1_2_port, B => n1349, Y => n4100)
                           ;
   U3961 : XNOR2X1 port map( A => results_b0_b1_4_port, B => n1347, Y => n4096)
                           ;
   U3962 : XNOR2X1 port map( A => results_b0_b1_6_port, B => n1345, Y => n4092)
                           ;
   U3963 : XNOR2X1 port map( A => results_b0_b1_8_port, B => n1343, Y => n4088)
                           ;
   U3964 : XNOR2X1 port map( A => results_b0_b1_10_port, B => n1358, Y => n4118
                           );
   U3965 : XNOR2X1 port map( A => results_b0_b1_12_port, B => n1356, Y => n4114
                           );
   U3966 : XNOR2X1 port map( A => results_b0_b1_14_port, B => n1354, Y => n4110
                           );
   U3967 : INVX1 port map( A => n169, Y => n1321);
   U3968 : INVX1 port map( A => n168, Y => n1341);
   U3969 : INVX1 port map( A => n166, Y => n1380);
   U3970 : INVX1 port map( A => n260, Y => n1238);
   U3971 : AOI32X1 port map( A0 => n1359, A1 => n4102, A2 => 
                           results_b0_b1_0_port, B0 => n1350, B1 => 
                           results_b0_b1_1_port, Y => n4101);
   U3972 : AOI22X1 port map( A0 => n1303, A1 => n1323, B0 => n4119, B1 => n4120
                           , Y => n4150);
   U3973 : AOI22X1 port map( A0 => n1318, A1 => n1338, B0 => n4148, B1 => n4149
                           , Y => n4146);
   U3974 : AOI22X1 port map( A0 => n1316, A1 => n1336, B0 => n4144, B1 => n4145
                           , Y => n4142);
   U3975 : XOR2X1 port map( A => n1320, B => n1340, Y => 
                           results_a1_a2_inv_0_port);
   U3976 : NOR2X1 port map( A => n220, B => n4545, Y => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b1);
   U3977 : NOR2X1 port map( A => n219, B => n4545, Y => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b2);
   U3978 : OAI2BB2X1 port map( B0 => n4122, B1 => n4121, A0N => n1304, A1N => 
                           n1324, Y => n4119);
   U3979 : OAI2BB2X1 port map( B0 => n4150, B1 => n4151, A0N => n1319, A1N => 
                           n1339, Y => n4148);
   U3980 : OAI2BB2X1 port map( B0 => n4146, B1 => n4147, A0N => n1317, A1N => 
                           n1337, Y => n4144);
   U3981 : OAI2BB2X1 port map( B0 => results_b0_b1_adderxn26, B1 => 
                           results_b0_b1_adderxn27, A0N => n1374, A1N => n1231,
                           Y => results_b0_b1_adderxn24);
   U3982 : OAI2BB2X1 port map( B0 => n4142, B1 => n4143, A0N => n1315, A1N => 
                           n1335, Y => n4140);
   U3983 : NOR2X1 port map( A => n220, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b1);
   U3984 : NOR2X1 port map( A => n220, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b1);
   U3985 : NOR2X1 port map( A => n220, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b1);
   U3986 : NOR2X1 port map( A => n219, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b2);
   U3987 : NOR2X1 port map( A => n219, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b2);
   U3988 : NOR2X1 port map( A => n219, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b2);
   U3989 : NOR2X1 port map( A => n218, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b3);
   U3990 : NOR2X1 port map( A => n218, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b3);
   U3991 : NOR2X1 port map( A => n217, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b4);
   U3992 : NOR2X1 port map( A => n217, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b4);
   U3993 : NOR2X1 port map( A => n216, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b5);
   U3994 : NOR2X1 port map( A => n216, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b5);
   U3995 : NOR2X1 port map( A => n216, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b5);
   U3996 : NOR2X1 port map( A => n215, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b6);
   U3997 : NOR2X1 port map( A => n215, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b6);
   U3998 : AOI22X1 port map( A0 => n4138, A1 => n1301, B0 => n1333, B1 => n1313
                           , Y => n4137);
   U3999 : NOR2X1 port map( A => n221, B => n4544, Y => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b0);
   U4000 : NOR2X1 port map( A => n231, B => n217, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b4);
   U4001 : NOR2X1 port map( A => n231, B => n218, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b3);
   U4002 : NOR2X1 port map( A => n231, B => n219, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b2);
   U4003 : NOR2X1 port map( A => n231, B => n215, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b6);
   U4004 : NOR2X1 port map( A => n221, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b0);
   U4005 : NOR2X1 port map( A => n219, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b2);
   U4006 : NOR2X1 port map( A => n219, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b2);
   U4007 : NOR2X1 port map( A => n218, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b3);
   U4008 : NOR2X1 port map( A => n218, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b3);
   U4009 : NOR2X1 port map( A => n217, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b4);
   U4010 : NOR2X1 port map( A => n217, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b4);
   U4011 : NOR2X1 port map( A => n216, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b5);
   U4012 : NOR2X1 port map( A => n216, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b5);
   U4013 : NOR2X1 port map( A => n215, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b6);
   U4014 : NOR2X1 port map( A => n215, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b6);
   U4015 : NOR2X1 port map( A => n222, B => n219, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b2);
   U4016 : NOR2X1 port map( A => n221, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b0);
   U4017 : NOR2X1 port map( A => n221, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b0);
   U4018 : NOR2X1 port map( A => n220, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b1);
   U4019 : NOR2X1 port map( A => n220, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b1);
   U4020 : NOR2X1 port map( A => n219, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b2);
   U4021 : NOR2X1 port map( A => n219, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b2);
   U4022 : NOR2X1 port map( A => n218, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b3);
   U4023 : NOR2X1 port map( A => n218, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b3);
   U4024 : NOR2X1 port map( A => n217, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b4);
   U4025 : NOR2X1 port map( A => n217, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b4);
   U4026 : NOR2X1 port map( A => n216, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b5);
   U4027 : NOR2X1 port map( A => n216, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b5);
   U4028 : NOR2X1 port map( A => n215, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b6);
   U4029 : NOR2X1 port map( A => n220, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b1);
   U4030 : NOR2X1 port map( A => n220, B => n225, Y => 
                           output_p1_times_a1_mul_componentxUMxa6_and_b1);
   U4031 : NOR2X1 port map( A => n221, B => n227, Y => 
                           output_p1_times_a1_mul_componentxUMxa4_and_b0);
   U4032 : NOR2X1 port map( A => n221, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b0);
   U4033 : XOR2X1 port map( A => n1359, B => results_b0_b1_0_port, Y => 
                           results_b0_b1_b2_0_port);
   U4034 : XOR2X1 port map( A => n1379, B => n1237, Y => results_b0_b1_0_port);
   U4035 : XOR2X1 port map( A => n1329, B => n1309, Y => n4132);
   U4036 : XOR2X1 port map( A => n1223, B => n1368, Y => 
                           results_b0_b1_adderxn15);
   U4037 : XOR2X1 port map( A => n1327, B => n1307, Y => n4128);
   U4038 : XOR2X1 port map( A => n1219, B => n1366, Y => 
                           results_b0_b1_adderxn11);
   U4039 : XOR2X1 port map( A => n1325, B => n1305, Y => n4124);
   U4040 : XOR2X1 port map( A => n1215, B => n1364, Y => results_b0_b1_adderxn7
                           );
   U4041 : XOR2X1 port map( A => n1323, B => n1303, Y => n4120);
   U4042 : XOR2X1 port map( A => n1211, B => n1362, Y => results_b0_b1_adderxn3
                           );
   U4043 : XOR2X1 port map( A => n1234, B => n1377, Y => 
                           results_b0_b1_adderxn33);
   U4044 : XOR2X1 port map( A => n1232, B => n1375, Y => 
                           results_b0_b1_adderxn29);
   U4045 : XOR2X1 port map( A => results_b0_b1_15_port, B => n1353, Y => n4108)
                           ;
   U4046 : XNOR2X1 port map( A => n100, B => n4135, Y => results_a1_a2_1_port);
   U4047 : NAND2X1 port map( A => n1340, B => n1320, Y => n100);
   U4048 : XOR2X1 port map( A => results_b0_b1_1_port, B => n1350, Y => n4102);
   U4049 : XNOR2X1 port map( A => n1330, B => n1310, Y => n4133);
   U4050 : XNOR2X1 port map( A => n1225, B => n1369, Y => 
                           results_b0_b1_adderxn16);
   U4051 : XNOR2X1 port map( A => n1328, B => n1308, Y => n4129);
   U4052 : XNOR2X1 port map( A => n1221, B => n1367, Y => 
                           results_b0_b1_adderxn12);
   U4053 : XNOR2X1 port map( A => n1326, B => n1306, Y => n4125);
   U4054 : XNOR2X1 port map( A => n1217, B => n1365, Y => 
                           results_b0_b1_adderxn8);
   U4055 : XNOR2X1 port map( A => n1324, B => n1304, Y => n4121);
   U4056 : XNOR2X1 port map( A => n1213, B => n1363, Y => 
                           results_b0_b1_adderxn4);
   U4057 : XNOR2X1 port map( A => n1235, B => n1378, Y => 
                           results_b0_b1_adderxn35);
   U4058 : XNOR2X1 port map( A => n1233, B => n1376, Y => 
                           results_b0_b1_adderxn31);
   U4059 : XNOR2X1 port map( A => n1231, B => n1374, Y => 
                           results_b0_b1_adderxn27);
   U4060 : XOR2X1 port map( A => results_b0_b1_16_port, B => n1352, Y => n4105)
                           ;
   U4061 : XNOR2X1 port map( A => n101, B => results_b0_b1_adderxn19, Y => 
                           results_b0_b1_1_port);
   U4062 : NAND2X1 port map( A => n1237, B => n1379, Y => n101);
   U4063 : XNOR2X1 port map( A => n102, B => n4102, Y => 
                           results_b0_b1_b2_1_port);
   U4064 : NAND2X1 port map( A => results_b0_b1_0_port, B => n1359, Y => n102);
   U4065 : XOR2X1 port map( A => results_a1_a2_inv_inverterxn10, B => 
                           results_a1_a2_17_port, Y => 
                           results_a1_a2_inv_17_port);
   U4066 : NAND2BX1 port map( AN => results_a1_a2_16_port, B => 
                           results_a1_a2_inv_inverterxn11, Y => 
                           results_a1_a2_inv_inverterxn10);
   U4067 : XOR2X1 port map( A => n4136, B => n4137, Y => results_a1_a2_17_port)
                           ;
   U4068 : XNOR2X1 port map( A => n1312, B => n1332, Y => n4136);
   U4069 : XOR2X1 port map( A => results_b0_b1_adderxn20, B => 
                           results_b0_b1_adderxn21, Y => results_b0_b1_17_port)
                           ;
   U4070 : XNOR2X1 port map( A => n1371, B => n1228, Y => 
                           results_b0_b1_adderxn20);
   U4071 : AOI22X1 port map( A0 => results_b0_b1_adderxn22, A1 => n1209, B0 => 
                           n1229, B1 => n1372, Y => results_b0_b1_adderxn21);
   U4072 : INVX1 port map( A => n4194, Y => n1371);
   U4073 : XOR2X1 port map( A => n4103, B => n4104, Y => 
                           results_b0_b1_b2_17_port);
   U4074 : XNOR2X1 port map( A => n1351, B => results_b0_b1_17_port, Y => n4103
                           );
   U4075 : AOI22X1 port map( A0 => n4105, A1 => n1207, B0 => 
                           results_b0_b1_16_port, B1 => n1352, Y => n4104);
   U4076 : INVX1 port map( A => n4250, Y => n1351);
   U4077 : INVX1 port map( A => n167, Y => n1360);
   U4078 : XNOR2X1 port map( A => n112, B => n360, Y => n4315);
   U4079 : INVX1 port map( A => results_b0_b1_adderxn23, Y => n1209);
   U4080 : AOI22X1 port map( A0 => n1373, A1 => n1230, B0 => 
                           results_b0_b1_adderxn24, B1 => 
                           results_b0_b1_adderxn25, Y => 
                           results_b0_b1_adderxn23);
   U4081 : INVX1 port map( A => n4139, Y => n1301);
   U4082 : AOI22X1 port map( A0 => n1314, A1 => n1334, B0 => n4140, B1 => n4141
                           , Y => n4139);
   U4083 : INVX1 port map( A => n4106, Y => n1207);
   U4084 : AOI22X1 port map( A0 => n1353, A1 => results_b0_b1_15_port, B0 => 
                           n4107, B1 => n4108, Y => n4106);
   U4085 : NOR2X1 port map( A => n218, B => n4545, Y => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b3);
   U4086 : NOR2X1 port map( A => n217, B => n4545, Y => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b4);
   U4087 : NOR2X1 port map( A => n220, B => n4542, Y => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b1);
   U4088 : NOR2X1 port map( A => n219, B => n4542, Y => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b2);
   U4089 : NOR2X1 port map( A => n215, B => n224, Y => 
                           output_p1_times_a1_mul_componentxUMxa7_and_b6);
   U4090 : NOR2X1 port map( A => n220, B => n4544, Y => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b1);
   U4091 : NOR2X1 port map( A => n219, B => n4544, Y => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b2);
   U4092 : NOR2X1 port map( A => n218, B => n4544, Y => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b3);
   U4093 : NOR2X1 port map( A => n221, B => n4543, Y => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b0);
   U4094 : NOR2X1 port map( A => n219, B => n4543, Y => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b2);
   U4095 : NOR2X1 port map( A => n220, B => n4543, Y => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b1);
   U4096 : NOR2X1 port map( A => n221, B => n4541, Y => 
                           output_p1_times_a1_mul_componentxUMxa14_and_b0);
   U4097 : NOR2X1 port map( A => n221, B => n228, Y => 
                           output_p1_times_a1_mul_componentxUMxa3_and_b0);
   U4098 : NOR2X1 port map( A => n221, B => n222, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b0);
   U4099 : NOR2X1 port map( A => n221, B => n229, Y => 
                           output_p1_times_a1_mul_componentxUMxa2_and_b0);
   U4100 : NOR2X1 port map( A => n222, B => n218, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b3);
   U4101 : NOR2X1 port map( A => n222, B => n217, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b4);
   U4102 : NOR2X1 port map( A => n220, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b1);
   U4103 : NOR2X1 port map( A => n222, B => n216, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b5);
   U4104 : NOR2X1 port map( A => n219, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b2);
   U4105 : NOR2X1 port map( A => n218, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b3);
   U4106 : NOR2X1 port map( A => n217, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b4);
   U4107 : NOR2X1 port map( A => n216, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b5);
   U4108 : NOR2X1 port map( A => n215, B => n226, Y => 
                           output_p1_times_a1_mul_componentxUMxa5_and_b6);
   U4109 : NOR2X1 port map( A => n215, B => n223, Y => 
                           output_p1_times_a1_mul_componentxUMxa8_and_b6);
   U4110 : NOR2X1 port map( A => n231, B => n220, Y => 
                           output_p1_times_a1_mul_componentxUMxa0_and_b1);
   U4111 : NOR2X1 port map( A => n222, B => n220, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b1);
   U4112 : NOR2X1 port map( A => n221, B => n4545, Y => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b0);
   U4113 : NOR2X1 port map( A => n221, B => n4542, Y => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b0);
   U4114 : NOR2X1 port map( A => n221, B => n230, Y => 
                           output_p1_times_a1_mul_componentxUMxa1_and_b0);
   U4115 : XOR2X1 port map( A => n1338, B => n1318, Y => n4149);
   U4116 : XOR2X1 port map( A => n1336, B => n1316, Y => n4145);
   U4117 : XOR2X1 port map( A => n1230, B => n1373, Y => 
                           results_b0_b1_adderxn25);
   U4118 : XOR2X1 port map( A => n1334, B => n1314, Y => n4141);
   U4119 : XNOR2X1 port map( A => n1339, B => n1319, Y => n4151);
   U4120 : XNOR2X1 port map( A => n1337, B => n1317, Y => n4147);
   U4121 : XNOR2X1 port map( A => n1335, B => n1315, Y => n4143);
   U4122 : XOR2X1 port map( A => n1229, B => n1372, Y => 
                           results_b0_b1_adderxn22);
   U4123 : XOR2X1 port map( A => n1333, B => n1313, Y => n4138);
   U4124 : NOR2X1 port map( A => n231, B => n221, Y => 
                           output_p1_times_a1_mul_componentxUMxfirst_vector_0_port);
   U4125 : NOR2X1 port map( A => n216, B => n4545, Y => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b5);
   U4126 : NOR2X1 port map( A => n215, B => n4545, Y => 
                           output_p1_times_a1_mul_componentxUMxa10_and_b6);
   U4127 : NOR2X1 port map( A => n218, B => n4542, Y => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b3);
   U4128 : NOR2X1 port map( A => n217, B => n4544, Y => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b4);
   U4129 : NOR2X1 port map( A => n216, B => n4544, Y => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b5);
   U4130 : NOR2X1 port map( A => n218, B => n4543, Y => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b3);
   U4131 : NOR2X1 port map( A => n217, B => n4543, Y => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b4);
   U4132 : NOR2X1 port map( A => n221, B => n4540, Y => 
                           output_p1_times_a1_mul_componentxUMxa15_and_b0);
   U4133 : NOR2X1 port map( A => n220, B => n4541, Y => 
                           output_p1_times_a1_mul_componentxUMxa14_and_b1);
   U4134 : NOR2X1 port map( A => n219, B => n4541, Y => 
                           output_p1_times_a1_mul_componentxUMxa14_and_b2);
   U4135 : NOR2X1 port map( A => n220, B => n4540, Y => 
                           output_p1_times_a1_mul_componentxUMxa15_and_b1);
   U4136 : NOR2X1 port map( A => n222, B => n215, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b6);
   U4137 : NOR2X1 port map( A => n217, B => n4542, Y => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b4);
   U4138 : NOR2X1 port map( A => n221, B => n4539, Y => 
                           output_p1_times_a1_mul_componentxUMxa16_and_b0);
   U4139 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa14_and_b3
                           , B => n3185, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715984_127849024_127850928);
   U4140 : NOR2X1 port map( A => n218, B => n4541, Y => 
                           output_p1_times_a1_mul_componentxUMxa14_and_b3);
   U4141 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa12_and_b5
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa13_and_b4, Y =>
                           n3185);
   U4142 : NOR2X1 port map( A => n216, B => n4543, Y => 
                           output_p1_times_a1_mul_componentxUMxa12_and_b5);
   U4143 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa15_and_b2
                           , B => 
                           output_p1_times_a1_mul_componentxUMxa16_and_b1, Y =>
                           n3186);
   U4144 : NOR2X1 port map( A => n219, B => n4540, Y => 
                           output_p1_times_a1_mul_componentxUMxa15_and_b2);
   U4145 : NOR2X1 port map( A => n220, B => n4539, Y => 
                           output_p1_times_a1_mul_componentxUMxa16_and_b1);
   U4146 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa11_and_b6
                           , B => n3184, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636480_127638384_127714080);
   U4147 : NOR2X1 port map( A => n215, B => n4544, Y => 
                           output_p1_times_a1_mul_componentxUMxa11_and_b6);
   U4148 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa9_and_b8,
                           B => output_p1_times_a1_mul_componentxUMxa10_and_b7,
                           Y => n3184);
   U4149 : NOR2X1 port map( A => n222, B => n213, Y => 
                           output_p1_times_a1_mul_componentxUMxa9_and_b8);
   U4150 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127627616_127629520_127824000, B 
                           => n3246, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer2_128199816_128200040_128199984);
   U4151 : XOR2X1 port map( A => output_p1_times_a1_mul_componentxUMxa17_and_b0
                           , B => n3186, Y => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127627616_127629520_127824000);
   U4152 : XOR2X1 port map( A => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127636480_127638384_127714080, B 
                           => 
                           output_p1_times_a1_mul_componentxUMxsum_layer1_127715984_127849024_127850928, Y 
                           => n3246);
   U4153 : NOR2X1 port map( A => n221, B => n9, Y => 
                           output_p1_times_a1_mul_componentxUMxa17_and_b0);
   U4154 : NOR2X1 port map( A => n178, B => n4439, Y => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b1);
   U4155 : NOR2X1 port map( A => n199, B => n4492, Y => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b1);
   U4156 : NOR2X1 port map( A => n241, B => n4598, Y => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b1);
   U4157 : NOR2X1 port map( A => n269, B => input_times_b0_mul_componentxn88, Y
                           => input_times_b0_mul_componentxUMxa10_and_b1);
   U4158 : NOR2X1 port map( A => n179, B => n4438, Y => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b0);
   U4159 : NOR2X1 port map( A => n270, B => input_times_b0_mul_componentxn87, Y
                           => input_times_b0_mul_componentxUMxa11_and_b0);
   U4160 : NOR2X1 port map( A => n180, B => n177, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b2);
   U4161 : NOR2X1 port map( A => n201, B => n198, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b2);
   U4162 : NOR2X1 port map( A => n243, B => n240, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b2);
   U4163 : NOR2X1 port map( A => n271, B => n268, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b2);
   U4164 : NOR2X1 port map( A => n177, B => n4439, Y => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b2);
   U4165 : NOR2X1 port map( A => n198, B => n4492, Y => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b2);
   U4166 : NOR2X1 port map( A => n240, B => n4598, Y => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b2);
   U4167 : NOR2X1 port map( A => n268, B => input_times_b0_mul_componentxn88, Y
                           => input_times_b0_mul_componentxUMxa10_and_b2);
   U4168 : NOR2X1 port map( A => n176, B => n4439, Y => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b3);
   U4169 : NOR2X1 port map( A => n197, B => n4492, Y => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b3);
   U4170 : NOR2X1 port map( A => n239, B => n4598, Y => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b3);
   U4171 : NOR2X1 port map( A => n267, B => input_times_b0_mul_componentxn88, Y
                           => input_times_b0_mul_componentxUMxa10_and_b3);
   U4172 : NOR2X1 port map( A => n175, B => n4439, Y => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b4);
   U4173 : NOR2X1 port map( A => n196, B => n4492, Y => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b4);
   U4174 : NOR2X1 port map( A => n238, B => n4598, Y => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b4);
   U4175 : NOR2X1 port map( A => n266, B => input_times_b0_mul_componentxn88, Y
                           => input_times_b0_mul_componentxUMxa10_and_b4);
   U4176 : NOR2X1 port map( A => n178, B => n4436, Y => 
                           input_p1_times_b1_mul_componentxUMxa13_and_b1);
   U4177 : NOR2X1 port map( A => n269, B => input_times_b0_mul_componentxn85, Y
                           => input_times_b0_mul_componentxUMxa13_and_b1);
   U4178 : NOR2X1 port map( A => n177, B => n4436, Y => 
                           input_p1_times_b1_mul_componentxUMxa13_and_b2);
   U4179 : NOR2X1 port map( A => n268, B => input_times_b0_mul_componentxn85, Y
                           => input_times_b0_mul_componentxUMxa13_and_b2);
   U4180 : NOR2X1 port map( A => n199, B => n4489, Y => 
                           input_p2_times_b2_mul_componentxUMxa13_and_b1);
   U4181 : NOR2X1 port map( A => n241, B => n4595, Y => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b1);
   U4182 : NOR2X1 port map( A => n198, B => n4489, Y => 
                           input_p2_times_b2_mul_componentxUMxa13_and_b2);
   U4183 : NOR2X1 port map( A => n240, B => n4595, Y => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b2);
   U4184 : NOR2X1 port map( A => n178, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b1);
   U4185 : NOR2X1 port map( A => n199, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b1);
   U4186 : NOR2X1 port map( A => n241, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b1);
   U4187 : NOR2X1 port map( A => n269, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b1);
   U4188 : NOR2X1 port map( A => n178, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b1);
   U4189 : NOR2X1 port map( A => n199, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b1);
   U4190 : NOR2X1 port map( A => n241, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b1);
   U4191 : NOR2X1 port map( A => n269, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b1);
   U4192 : NOR2X1 port map( A => n177, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b2);
   U4193 : NOR2X1 port map( A => n198, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b2);
   U4194 : NOR2X1 port map( A => n240, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b2);
   U4195 : NOR2X1 port map( A => n268, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b2);
   U4196 : NOR2X1 port map( A => n177, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b2);
   U4197 : NOR2X1 port map( A => n198, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b2);
   U4198 : NOR2X1 port map( A => n240, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b2);
   U4199 : NOR2X1 port map( A => n268, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b2);
   U4200 : NOR2X1 port map( A => n177, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b2);
   U4201 : NOR2X1 port map( A => n198, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b2);
   U4202 : NOR2X1 port map( A => n240, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b2);
   U4203 : NOR2X1 port map( A => n268, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b2);
   U4204 : NOR2X1 port map( A => n176, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b3);
   U4205 : NOR2X1 port map( A => n197, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b3);
   U4206 : NOR2X1 port map( A => n239, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b3);
   U4207 : NOR2X1 port map( A => n267, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b3);
   U4208 : NOR2X1 port map( A => n176, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b3);
   U4209 : NOR2X1 port map( A => n197, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b3);
   U4210 : NOR2X1 port map( A => n239, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b3);
   U4211 : NOR2X1 port map( A => n267, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b3);
   U4212 : NOR2X1 port map( A => n176, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b3);
   U4213 : NOR2X1 port map( A => n197, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b3);
   U4214 : NOR2X1 port map( A => n239, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b3);
   U4215 : NOR2X1 port map( A => n267, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b3);
   U4216 : NOR2X1 port map( A => n175, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b4);
   U4217 : NOR2X1 port map( A => n196, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b4);
   U4218 : NOR2X1 port map( A => n238, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b4);
   U4219 : NOR2X1 port map( A => n266, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b4);
   U4220 : NOR2X1 port map( A => n175, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b4);
   U4221 : NOR2X1 port map( A => n196, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b4);
   U4222 : NOR2X1 port map( A => n238, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b4);
   U4223 : NOR2X1 port map( A => n266, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b4);
   U4224 : NOR2X1 port map( A => n175, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b4);
   U4225 : NOR2X1 port map( A => n196, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b4);
   U4226 : NOR2X1 port map( A => n238, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b4);
   U4227 : NOR2X1 port map( A => n266, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b4);
   U4228 : NOR2X1 port map( A => n174, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b5);
   U4229 : NOR2X1 port map( A => n195, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b5);
   U4230 : NOR2X1 port map( A => n237, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b5);
   U4231 : NOR2X1 port map( A => n265, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b5);
   U4232 : NOR2X1 port map( A => n174, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b5);
   U4233 : NOR2X1 port map( A => n195, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b5);
   U4234 : NOR2X1 port map( A => n237, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b5);
   U4235 : NOR2X1 port map( A => n265, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b5);
   U4236 : NOR2X1 port map( A => n174, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b5);
   U4237 : NOR2X1 port map( A => n195, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b5);
   U4238 : NOR2X1 port map( A => n237, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b5);
   U4239 : NOR2X1 port map( A => n265, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b5);
   U4240 : NOR2X1 port map( A => n172, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b7);
   U4241 : NOR2X1 port map( A => n173, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b6);
   U4242 : NOR2X1 port map( A => n194, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b6);
   U4243 : NOR2X1 port map( A => n236, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b6);
   U4244 : NOR2X1 port map( A => n263, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b7);
   U4245 : NOR2X1 port map( A => n264, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b6);
   U4246 : NOR2X1 port map( A => n173, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b6);
   U4247 : NOR2X1 port map( A => n194, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b6);
   U4248 : NOR2X1 port map( A => n236, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b6);
   U4249 : NOR2X1 port map( A => n264, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b6);
   U4250 : NOR2X1 port map( A => n193, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b7);
   U4251 : NOR2X1 port map( A => n235, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b7);
   U4252 : NOR2X1 port map( A => n172, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b7);
   U4253 : NOR2X1 port map( A => n263, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b7);
   U4254 : NOR2X1 port map( A => n178, B => n4438, Y => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b1);
   U4255 : NOR2X1 port map( A => n269, B => input_times_b0_mul_componentxn87, Y
                           => input_times_b0_mul_componentxUMxa11_and_b1);
   U4256 : NOR2X1 port map( A => n177, B => n4438, Y => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b2);
   U4257 : NOR2X1 port map( A => n268, B => input_times_b0_mul_componentxn87, Y
                           => input_times_b0_mul_componentxUMxa11_and_b2);
   U4258 : NOR2X1 port map( A => n176, B => n4438, Y => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b3);
   U4259 : NOR2X1 port map( A => n267, B => input_times_b0_mul_componentxn87, Y
                           => input_times_b0_mul_componentxUMxa11_and_b3);
   U4260 : NOR2X1 port map( A => n179, B => n4437, Y => 
                           input_p1_times_b1_mul_componentxUMxa12_and_b0);
   U4261 : NOR2X1 port map( A => n270, B => input_times_b0_mul_componentxn86, Y
                           => input_times_b0_mul_componentxUMxa12_and_b0);
   U4262 : NOR2X1 port map( A => n177, B => n4437, Y => 
                           input_p1_times_b1_mul_componentxUMxa12_and_b2);
   U4263 : NOR2X1 port map( A => n268, B => input_times_b0_mul_componentxn86, Y
                           => input_times_b0_mul_componentxUMxa12_and_b2);
   U4264 : NOR2X1 port map( A => n200, B => n4491, Y => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b0);
   U4265 : NOR2X1 port map( A => n242, B => n4597, Y => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b0);
   U4266 : NOR2X1 port map( A => n199, B => n4491, Y => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b1);
   U4267 : NOR2X1 port map( A => n241, B => n4597, Y => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b1);
   U4268 : NOR2X1 port map( A => n198, B => n4491, Y => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b2);
   U4269 : NOR2X1 port map( A => n240, B => n4597, Y => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b2);
   U4270 : NOR2X1 port map( A => n197, B => n4491, Y => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b3);
   U4271 : NOR2X1 port map( A => n239, B => n4597, Y => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b3);
   U4272 : NOR2X1 port map( A => n200, B => n4490, Y => 
                           input_p2_times_b2_mul_componentxUMxa12_and_b0);
   U4273 : NOR2X1 port map( A => n242, B => n4596, Y => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b0);
   U4274 : NOR2X1 port map( A => n198, B => n4490, Y => 
                           input_p2_times_b2_mul_componentxUMxa12_and_b2);
   U4275 : NOR2X1 port map( A => n240, B => n4596, Y => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b2);
   U4276 : NOR2X1 port map( A => n179, B => n4434, Y => 
                           input_p1_times_b1_mul_componentxUMxa15_and_b0);
   U4277 : NOR2X1 port map( A => n270, B => input_times_b0_mul_componentxn83, Y
                           => input_times_b0_mul_componentxUMxa15_and_b0);
   U4278 : NOR2X1 port map( A => n179, B => n4435, Y => 
                           input_p1_times_b1_mul_componentxUMxa14_and_b0);
   U4279 : NOR2X1 port map( A => n270, B => input_times_b0_mul_componentxn84, Y
                           => input_times_b0_mul_componentxUMxa14_and_b0);
   U4280 : NOR2X1 port map( A => n178, B => n4437, Y => 
                           input_p1_times_b1_mul_componentxUMxa12_and_b1);
   U4281 : NOR2X1 port map( A => n269, B => input_times_b0_mul_componentxn86, Y
                           => input_times_b0_mul_componentxUMxa12_and_b1);
   U4282 : NOR2X1 port map( A => n200, B => n4487, Y => 
                           input_p2_times_b2_mul_componentxUMxa15_and_b0);
   U4283 : NOR2X1 port map( A => n242, B => n4593, Y => 
                           output_p2_times_a2_mul_componentxUMxa15_and_b0);
   U4284 : NOR2X1 port map( A => n199, B => n4490, Y => 
                           input_p2_times_b2_mul_componentxUMxa12_and_b1);
   U4285 : NOR2X1 port map( A => n241, B => n4596, Y => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b1);
   U4286 : NOR2X1 port map( A => n200, B => n4488, Y => 
                           input_p2_times_b2_mul_componentxUMxa14_and_b0);
   U4287 : NOR2X1 port map( A => n242, B => n4594, Y => 
                           output_p2_times_a2_mul_componentxUMxa14_and_b0);
   U4288 : NOR2X1 port map( A => n189, B => n175, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b4);
   U4289 : NOR2X1 port map( A => n280, B => n266, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b4);
   U4290 : NOR2X1 port map( A => n189, B => n174, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b5);
   U4291 : NOR2X1 port map( A => n280, B => n265, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b5);
   U4292 : NOR2X1 port map( A => n189, B => n176, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b3);
   U4293 : NOR2X1 port map( A => n280, B => n267, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b3);
   U4294 : NOR2X1 port map( A => n189, B => n171, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b8);
   U4295 : NOR2X1 port map( A => n189, B => n172, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b7);
   U4296 : NOR2X1 port map( A => n280, B => n262, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b8);
   U4297 : NOR2X1 port map( A => n280, B => n263, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b7);
   U4298 : NOR2X1 port map( A => n189, B => n173, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b6);
   U4299 : NOR2X1 port map( A => n280, B => n264, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b6);
   U4300 : NOR2X1 port map( A => n210, B => n196, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b4);
   U4301 : NOR2X1 port map( A => n252, B => n238, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b4);
   U4302 : NOR2X1 port map( A => n210, B => n195, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b5);
   U4303 : NOR2X1 port map( A => n252, B => n237, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b5);
   U4304 : NOR2X1 port map( A => n210, B => n197, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b3);
   U4305 : NOR2X1 port map( A => n252, B => n239, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b3);
   U4306 : NOR2X1 port map( A => n210, B => n192, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b8);
   U4307 : NOR2X1 port map( A => n210, B => n193, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b7);
   U4308 : NOR2X1 port map( A => n252, B => n234, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b8);
   U4309 : NOR2X1 port map( A => n252, B => n235, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b7);
   U4310 : NOR2X1 port map( A => n210, B => n194, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b6);
   U4311 : NOR2X1 port map( A => n252, B => n236, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b6);
   U4312 : NOR2X1 port map( A => n179, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b0);
   U4313 : NOR2X1 port map( A => n200, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b0);
   U4314 : NOR2X1 port map( A => n242, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b0);
   U4315 : NOR2X1 port map( A => n270, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b0);
   U4316 : NOR2X1 port map( A => n179, B => n180, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b0);
   U4317 : NOR2X1 port map( A => n200, B => n201, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b0);
   U4318 : NOR2X1 port map( A => n242, B => n243, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b0);
   U4319 : NOR2X1 port map( A => n270, B => n271, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b0);
   U4320 : NOR2X1 port map( A => n177, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b2);
   U4321 : NOR2X1 port map( A => n198, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b2);
   U4322 : NOR2X1 port map( A => n240, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b2);
   U4323 : NOR2X1 port map( A => n268, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b2);
   U4324 : NOR2X1 port map( A => n177, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b2);
   U4325 : NOR2X1 port map( A => n198, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b2);
   U4326 : NOR2X1 port map( A => n240, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b2);
   U4327 : NOR2X1 port map( A => n268, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b2);
   U4328 : NOR2X1 port map( A => n176, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b3);
   U4329 : NOR2X1 port map( A => n197, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b3);
   U4330 : NOR2X1 port map( A => n239, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b3);
   U4331 : NOR2X1 port map( A => n267, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b3);
   U4332 : NOR2X1 port map( A => n176, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b3);
   U4333 : NOR2X1 port map( A => n197, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b3);
   U4334 : NOR2X1 port map( A => n239, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b3);
   U4335 : NOR2X1 port map( A => n267, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b3);
   U4336 : NOR2X1 port map( A => n175, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b4);
   U4337 : NOR2X1 port map( A => n196, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b4);
   U4338 : NOR2X1 port map( A => n238, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b4);
   U4339 : NOR2X1 port map( A => n266, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b4);
   U4340 : NOR2X1 port map( A => n175, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b4);
   U4341 : NOR2X1 port map( A => n196, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b4);
   U4342 : NOR2X1 port map( A => n238, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b4);
   U4343 : NOR2X1 port map( A => n266, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b4);
   U4344 : NOR2X1 port map( A => n174, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b5);
   U4345 : NOR2X1 port map( A => n195, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b5);
   U4346 : NOR2X1 port map( A => n237, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b5);
   U4347 : NOR2X1 port map( A => n265, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b5);
   U4348 : NOR2X1 port map( A => n174, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b5);
   U4349 : NOR2X1 port map( A => n195, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b5);
   U4350 : NOR2X1 port map( A => n237, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b5);
   U4351 : NOR2X1 port map( A => n265, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b5);
   U4352 : NOR2X1 port map( A => n173, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b6);
   U4353 : NOR2X1 port map( A => n264, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b6);
   U4354 : NOR2X1 port map( A => n173, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b6);
   U4355 : NOR2X1 port map( A => n194, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b6);
   U4356 : NOR2X1 port map( A => n236, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b6);
   U4357 : NOR2X1 port map( A => n264, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b6);
   U4358 : NOR2X1 port map( A => n179, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b0);
   U4359 : NOR2X1 port map( A => n200, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b0);
   U4360 : NOR2X1 port map( A => n242, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b0);
   U4361 : NOR2X1 port map( A => n270, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b0);
   U4362 : NOR2X1 port map( A => n179, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b0);
   U4363 : NOR2X1 port map( A => n200, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b0);
   U4364 : NOR2X1 port map( A => n242, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b0);
   U4365 : NOR2X1 port map( A => n270, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b0);
   U4366 : NOR2X1 port map( A => n180, B => n176, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b3);
   U4367 : NOR2X1 port map( A => n201, B => n197, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b3);
   U4368 : NOR2X1 port map( A => n243, B => n239, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b3);
   U4369 : NOR2X1 port map( A => n271, B => n267, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b3);
   U4370 : NOR2X1 port map( A => n172, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b7);
   U4371 : NOR2X1 port map( A => n193, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b7);
   U4372 : NOR2X1 port map( A => n235, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b7);
   U4373 : NOR2X1 port map( A => n263, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b7);
   U4374 : NOR2X1 port map( A => n180, B => n175, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b4);
   U4375 : NOR2X1 port map( A => n201, B => n196, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b4);
   U4376 : NOR2X1 port map( A => n243, B => n238, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b4);
   U4377 : NOR2X1 port map( A => n271, B => n266, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b4);
   U4378 : NOR2X1 port map( A => n178, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b1);
   U4379 : NOR2X1 port map( A => n199, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b1);
   U4380 : NOR2X1 port map( A => n241, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b1);
   U4381 : NOR2X1 port map( A => n269, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b1);
   U4382 : NOR2X1 port map( A => n178, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b1);
   U4383 : NOR2X1 port map( A => n199, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b1);
   U4384 : NOR2X1 port map( A => n241, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b1);
   U4385 : NOR2X1 port map( A => n269, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b1);
   U4386 : NOR2X1 port map( A => n180, B => n174, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b5);
   U4387 : NOR2X1 port map( A => n201, B => n195, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b5);
   U4388 : NOR2X1 port map( A => n243, B => n237, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b5);
   U4389 : NOR2X1 port map( A => n271, B => n265, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b5);
   U4390 : NOR2X1 port map( A => n177, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b2);
   U4391 : NOR2X1 port map( A => n198, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b2);
   U4392 : NOR2X1 port map( A => n240, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b2);
   U4393 : NOR2X1 port map( A => n268, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b2);
   U4394 : NOR2X1 port map( A => n177, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b2);
   U4395 : NOR2X1 port map( A => n198, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b2);
   U4396 : NOR2X1 port map( A => n240, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b2);
   U4397 : NOR2X1 port map( A => n268, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b2);
   U4398 : NOR2X1 port map( A => n177, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b2);
   U4399 : NOR2X1 port map( A => n198, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b2);
   U4400 : NOR2X1 port map( A => n240, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b2);
   U4401 : NOR2X1 port map( A => n268, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b2);
   U4402 : NOR2X1 port map( A => n176, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b3);
   U4403 : NOR2X1 port map( A => n197, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b3);
   U4404 : NOR2X1 port map( A => n239, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b3);
   U4405 : NOR2X1 port map( A => n267, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b3);
   U4406 : NOR2X1 port map( A => n176, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b3);
   U4407 : NOR2X1 port map( A => n197, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b3);
   U4408 : NOR2X1 port map( A => n239, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b3);
   U4409 : NOR2X1 port map( A => n267, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b3);
   U4410 : NOR2X1 port map( A => n176, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b3);
   U4411 : NOR2X1 port map( A => n197, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b3);
   U4412 : NOR2X1 port map( A => n239, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b3);
   U4413 : NOR2X1 port map( A => n267, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b3);
   U4414 : NOR2X1 port map( A => n175, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b4);
   U4415 : NOR2X1 port map( A => n196, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b4);
   U4416 : NOR2X1 port map( A => n238, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b4);
   U4417 : NOR2X1 port map( A => n266, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b4);
   U4418 : NOR2X1 port map( A => n175, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b4);
   U4419 : NOR2X1 port map( A => n196, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b4);
   U4420 : NOR2X1 port map( A => n238, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b4);
   U4421 : NOR2X1 port map( A => n266, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b4);
   U4422 : NOR2X1 port map( A => n174, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b5);
   U4423 : NOR2X1 port map( A => n195, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b5);
   U4424 : NOR2X1 port map( A => n237, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b5);
   U4425 : NOR2X1 port map( A => n265, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b5);
   U4426 : NOR2X1 port map( A => n174, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b5);
   U4427 : NOR2X1 port map( A => n265, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b5);
   U4428 : NOR2X1 port map( A => n178, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b1);
   U4429 : NOR2X1 port map( A => n199, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b1);
   U4430 : NOR2X1 port map( A => n241, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b1);
   U4431 : NOR2X1 port map( A => n269, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b1);
   U4432 : NOR2X1 port map( A => n178, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b1);
   U4433 : NOR2X1 port map( A => n199, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b1);
   U4434 : NOR2X1 port map( A => n241, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b1);
   U4435 : NOR2X1 port map( A => n269, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b1);
   U4436 : NOR2X1 port map( A => n180, B => n178, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b1);
   U4437 : NOR2X1 port map( A => n201, B => n199, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b1);
   U4438 : NOR2X1 port map( A => n243, B => n241, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b1);
   U4439 : NOR2X1 port map( A => n271, B => n269, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b1);
   U4440 : NOR2X1 port map( A => n179, B => n4439, Y => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b0);
   U4441 : NOR2X1 port map( A => n200, B => n4492, Y => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b0);
   U4442 : NOR2X1 port map( A => n242, B => n4598, Y => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b0);
   U4443 : NOR2X1 port map( A => n270, B => input_times_b0_mul_componentxn88, Y
                           => input_times_b0_mul_componentxUMxa10_and_b0);
   U4444 : NOR2X1 port map( A => n179, B => n4436, Y => 
                           input_p1_times_b1_mul_componentxUMxa13_and_b0);
   U4445 : NOR2X1 port map( A => n270, B => input_times_b0_mul_componentxn85, Y
                           => input_times_b0_mul_componentxUMxa13_and_b0);
   U4446 : NOR2X1 port map( A => n200, B => n4489, Y => 
                           input_p2_times_b2_mul_componentxUMxa13_and_b0);
   U4447 : NOR2X1 port map( A => n242, B => n4595, Y => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b0);
   U4448 : NOR2X1 port map( A => n179, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b0);
   U4449 : NOR2X1 port map( A => n200, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b0);
   U4450 : NOR2X1 port map( A => n242, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b0);
   U4451 : NOR2X1 port map( A => n270, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b0);
   U4452 : NOR2X1 port map( A => n179, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b0);
   U4453 : NOR2X1 port map( A => n200, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b0);
   U4454 : NOR2X1 port map( A => n242, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b0);
   U4455 : NOR2X1 port map( A => n270, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b0);
   U4456 : NOR2X1 port map( A => n4422, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b10);
   U4457 : NOR2X1 port map( A => n4475, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b10);
   U4458 : NOR2X1 port map( A => n4581, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b10);
   U4459 : NOR2X1 port map( A => input_times_b0_mul_componentxn71, B => n279, Y
                           => input_times_b0_mul_componentxUMxa1_and_b10);
   U4460 : NOR2X1 port map( A => n4422, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b10);
   U4461 : NOR2X1 port map( A => n4475, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b10);
   U4462 : NOR2X1 port map( A => n4581, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b10);
   U4463 : NOR2X1 port map( A => input_times_b0_mul_componentxn71, B => n276, Y
                           => input_times_b0_mul_componentxUMxa4_and_b10);
   U4464 : NOR2X1 port map( A => n174, B => n4439, Y => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b5);
   U4465 : NOR2X1 port map( A => n195, B => n4492, Y => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b5);
   U4466 : NOR2X1 port map( A => n237, B => n4598, Y => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b5);
   U4467 : NOR2X1 port map( A => n265, B => input_times_b0_mul_componentxn88, Y
                           => input_times_b0_mul_componentxUMxa10_and_b5);
   U4468 : NOR2X1 port map( A => n173, B => n4439, Y => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b6);
   U4469 : NOR2X1 port map( A => n194, B => n4492, Y => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b6);
   U4470 : NOR2X1 port map( A => n236, B => n4598, Y => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b6);
   U4471 : NOR2X1 port map( A => n264, B => input_times_b0_mul_componentxn88, Y
                           => input_times_b0_mul_componentxUMxa10_and_b6);
   U4472 : NOR2X1 port map( A => n4421, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b11);
   U4473 : NOR2X1 port map( A => n4474, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b11);
   U4474 : NOR2X1 port map( A => n4580, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b11);
   U4475 : NOR2X1 port map( A => input_times_b0_mul_componentxn70, B => n279, Y
                           => input_times_b0_mul_componentxUMxa1_and_b11);
   U4476 : NOR2X1 port map( A => n4420, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b12);
   U4477 : NOR2X1 port map( A => n4473, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b12);
   U4478 : NOR2X1 port map( A => n4579, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b12);
   U4479 : NOR2X1 port map( A => input_times_b0_mul_componentxn69, B => n279, Y
                           => input_times_b0_mul_componentxUMxa1_and_b12);
   U4480 : NOR2X1 port map( A => n176, B => n4436, Y => 
                           input_p1_times_b1_mul_componentxUMxa13_and_b3);
   U4481 : NOR2X1 port map( A => n267, B => input_times_b0_mul_componentxn85, Y
                           => input_times_b0_mul_componentxUMxa13_and_b3);
   U4482 : NOR2X1 port map( A => n197, B => n4489, Y => 
                           input_p2_times_b2_mul_componentxUMxa13_and_b3);
   U4483 : NOR2X1 port map( A => n239, B => n4595, Y => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b3);
   U4484 : NOR2X1 port map( A => n178, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b1);
   U4485 : NOR2X1 port map( A => n199, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b1);
   U4486 : NOR2X1 port map( A => n241, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b1);
   U4487 : NOR2X1 port map( A => n269, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b1);
   U4488 : NOR2X1 port map( A => n171, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b8);
   U4489 : NOR2X1 port map( A => n262, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b8);
   U4490 : NOR2X1 port map( A => n170, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b9);
   U4491 : NOR2X1 port map( A => n261, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b9);
   U4492 : NOR2X1 port map( A => n173, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b6);
   U4493 : NOR2X1 port map( A => n194, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b6);
   U4494 : NOR2X1 port map( A => n236, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b6);
   U4495 : NOR2X1 port map( A => n264, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b6);
   U4496 : NOR2X1 port map( A => n192, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b8);
   U4497 : NOR2X1 port map( A => n234, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b8);
   U4498 : NOR2X1 port map( A => n191, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b9);
   U4499 : NOR2X1 port map( A => n233, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b9);
   U4500 : NOR2X1 port map( A => n172, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b7);
   U4501 : NOR2X1 port map( A => n193, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b7);
   U4502 : NOR2X1 port map( A => n235, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b7);
   U4503 : NOR2X1 port map( A => n263, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b7);
   U4504 : NOR2X1 port map( A => n193, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b7);
   U4505 : NOR2X1 port map( A => n235, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b7);
   U4506 : NOR2X1 port map( A => n171, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b8);
   U4507 : NOR2X1 port map( A => n262, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b8);
   U4508 : NOR2X1 port map( A => n170, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b9);
   U4509 : NOR2X1 port map( A => n261, B => n276, Y => 
                           input_times_b0_mul_componentxUMxa4_and_b9);
   U4510 : NOR2X1 port map( A => n192, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b8);
   U4511 : NOR2X1 port map( A => n234, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b8);
   U4512 : NOR2X1 port map( A => n191, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b9);
   U4513 : NOR2X1 port map( A => n233, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b9);
   U4514 : NOR2X1 port map( A => n171, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b8);
   U4515 : NOR2X1 port map( A => n262, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b8);
   U4516 : NOR2X1 port map( A => n4422, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b10);
   U4517 : NOR2X1 port map( A => n4475, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b10);
   U4518 : NOR2X1 port map( A => n4581, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b10);
   U4519 : NOR2X1 port map( A => input_times_b0_mul_componentxn71, B => n277, Y
                           => input_times_b0_mul_componentxUMxa3_and_b10);
   U4520 : NOR2X1 port map( A => n189, B => n4422, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b10);
   U4521 : NOR2X1 port map( A => n210, B => n4475, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b10);
   U4522 : NOR2X1 port map( A => n252, B => n4581, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b10);
   U4523 : NOR2X1 port map( A => n280, B => input_times_b0_mul_componentxn71, Y
                           => input_times_b0_mul_componentxUMxa0_and_b10);
   U4524 : NOR2X1 port map( A => n4422, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b10);
   U4525 : NOR2X1 port map( A => n4475, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b10);
   U4526 : NOR2X1 port map( A => n4581, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b10);
   U4527 : NOR2X1 port map( A => input_times_b0_mul_componentxn71, B => n278, Y
                           => input_times_b0_mul_componentxUMxa2_and_b10);
   U4528 : NOR2X1 port map( A => n4421, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b11);
   U4529 : NOR2X1 port map( A => n4474, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b11);
   U4530 : NOR2X1 port map( A => n4580, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b11);
   U4531 : NOR2X1 port map( A => input_times_b0_mul_componentxn70, B => n277, Y
                           => input_times_b0_mul_componentxUMxa3_and_b11);
   U4532 : NOR2X1 port map( A => n189, B => n4421, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b11);
   U4533 : NOR2X1 port map( A => n210, B => n4474, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b11);
   U4534 : NOR2X1 port map( A => n252, B => n4580, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b11);
   U4535 : NOR2X1 port map( A => n280, B => input_times_b0_mul_componentxn70, Y
                           => input_times_b0_mul_componentxUMxa0_and_b11);
   U4536 : NOR2X1 port map( A => n4421, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b11);
   U4537 : NOR2X1 port map( A => n4474, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b11);
   U4538 : NOR2X1 port map( A => n4580, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b11);
   U4539 : NOR2X1 port map( A => input_times_b0_mul_componentxn70, B => n278, Y
                           => input_times_b0_mul_componentxUMxa2_and_b11);
   U4540 : NOR2X1 port map( A => n175, B => n4438, Y => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b4);
   U4541 : NOR2X1 port map( A => n266, B => input_times_b0_mul_componentxn87, Y
                           => input_times_b0_mul_componentxUMxa11_and_b4);
   U4542 : NOR2X1 port map( A => n174, B => n4438, Y => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b5);
   U4543 : NOR2X1 port map( A => n265, B => input_times_b0_mul_componentxn87, Y
                           => input_times_b0_mul_componentxUMxa11_and_b5);
   U4544 : NOR2X1 port map( A => n176, B => n4437, Y => 
                           input_p1_times_b1_mul_componentxUMxa12_and_b3);
   U4545 : NOR2X1 port map( A => n267, B => input_times_b0_mul_componentxn86, Y
                           => input_times_b0_mul_componentxUMxa12_and_b3);
   U4546 : NOR2X1 port map( A => n175, B => n4437, Y => 
                           input_p1_times_b1_mul_componentxUMxa12_and_b4);
   U4547 : NOR2X1 port map( A => n266, B => input_times_b0_mul_componentxn86, Y
                           => input_times_b0_mul_componentxUMxa12_and_b4);
   U4548 : NOR2X1 port map( A => n189, B => n4420, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b12);
   U4549 : NOR2X1 port map( A => n210, B => n4473, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b12);
   U4550 : NOR2X1 port map( A => n252, B => n4579, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b12);
   U4551 : NOR2X1 port map( A => n280, B => input_times_b0_mul_componentxn69, Y
                           => input_times_b0_mul_componentxUMxa0_and_b12);
   U4552 : NOR2X1 port map( A => n196, B => n4491, Y => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b4);
   U4553 : NOR2X1 port map( A => n238, B => n4597, Y => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b4);
   U4554 : NOR2X1 port map( A => n195, B => n4491, Y => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b5);
   U4555 : NOR2X1 port map( A => n237, B => n4597, Y => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b5);
   U4556 : NOR2X1 port map( A => n197, B => n4490, Y => 
                           input_p2_times_b2_mul_componentxUMxa12_and_b3);
   U4557 : NOR2X1 port map( A => n239, B => n4596, Y => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b3);
   U4558 : NOR2X1 port map( A => n196, B => n4490, Y => 
                           input_p2_times_b2_mul_componentxUMxa12_and_b4);
   U4559 : NOR2X1 port map( A => n238, B => n4596, Y => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b4);
   U4560 : NOR2X1 port map( A => n280, B => input_times_b0_mul_componentxn68, Y
                           => input_times_b0_mul_componentxUMxa0_and_b13);
   U4561 : NOR2X1 port map( A => n189, B => n4419, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b13);
   U4562 : NOR2X1 port map( A => n210, B => n4472, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b13);
   U4563 : NOR2X1 port map( A => n252, B => n4578, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b13);
   U4564 : NOR2X1 port map( A => n178, B => n4435, Y => 
                           input_p1_times_b1_mul_componentxUMxa14_and_b1);
   U4565 : NOR2X1 port map( A => n269, B => input_times_b0_mul_componentxn84, Y
                           => input_times_b0_mul_componentxUMxa14_and_b1);
   U4566 : NOR2X1 port map( A => n177, B => n4435, Y => 
                           input_p1_times_b1_mul_componentxUMxa14_and_b2);
   U4567 : NOR2X1 port map( A => n268, B => input_times_b0_mul_componentxn84, Y
                           => input_times_b0_mul_componentxUMxa14_and_b2);
   U4568 : NOR2X1 port map( A => n199, B => n4488, Y => 
                           input_p2_times_b2_mul_componentxUMxa14_and_b1);
   U4569 : NOR2X1 port map( A => n241, B => n4594, Y => 
                           output_p2_times_a2_mul_componentxUMxa14_and_b1);
   U4570 : NOR2X1 port map( A => n198, B => n4488, Y => 
                           input_p2_times_b2_mul_componentxUMxa14_and_b2);
   U4571 : NOR2X1 port map( A => n240, B => n4594, Y => 
                           output_p2_times_a2_mul_componentxUMxa14_and_b2);
   U4572 : NOR2X1 port map( A => n178, B => n4434, Y => 
                           input_p1_times_b1_mul_componentxUMxa15_and_b1);
   U4573 : NOR2X1 port map( A => n269, B => input_times_b0_mul_componentxn83, Y
                           => input_times_b0_mul_componentxUMxa15_and_b1);
   U4574 : NOR2X1 port map( A => n189, B => n177, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b2);
   U4575 : NOR2X1 port map( A => n280, B => n268, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b2);
   U4576 : NOR2X1 port map( A => n189, B => n170, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b9);
   U4577 : NOR2X1 port map( A => n280, B => n261, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b9);
   U4578 : NOR2X1 port map( A => n210, B => n198, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b2);
   U4579 : NOR2X1 port map( A => n252, B => n240, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b2);
   U4580 : NOR2X1 port map( A => n210, B => n191, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b9);
   U4581 : NOR2X1 port map( A => n252, B => n233, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b9);
   U4582 : NOR2X1 port map( A => n179, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b0);
   U4583 : NOR2X1 port map( A => n200, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b0);
   U4584 : NOR2X1 port map( A => n242, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b0);
   U4585 : NOR2X1 port map( A => n270, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b0);
   U4586 : NOR2X1 port map( A => n199, B => n4487, Y => 
                           input_p2_times_b2_mul_componentxUMxa15_and_b1);
   U4587 : NOR2X1 port map( A => n241, B => n4593, Y => 
                           output_p2_times_a2_mul_componentxUMxa15_and_b1);
   U4588 : NOR2X1 port map( A => n194, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b6);
   U4589 : NOR2X1 port map( A => n236, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b6);
   U4590 : NOR2X1 port map( A => n179, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b0);
   U4591 : NOR2X1 port map( A => n200, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b0);
   U4592 : NOR2X1 port map( A => n242, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b0);
   U4593 : NOR2X1 port map( A => n270, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b0);
   U4594 : NOR2X1 port map( A => n172, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b7);
   U4595 : NOR2X1 port map( A => n193, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b7);
   U4596 : NOR2X1 port map( A => n235, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b7);
   U4597 : NOR2X1 port map( A => n263, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b7);
   U4598 : NOR2X1 port map( A => n170, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b9);
   U4599 : NOR2X1 port map( A => n261, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b9);
   U4600 : NOR2X1 port map( A => n171, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b8);
   U4601 : NOR2X1 port map( A => n262, B => n277, Y => 
                           input_times_b0_mul_componentxUMxa3_and_b8);
   U4602 : NOR2X1 port map( A => n191, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b9);
   U4603 : NOR2X1 port map( A => n233, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b9);
   U4604 : NOR2X1 port map( A => n192, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b8);
   U4605 : NOR2X1 port map( A => n234, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b8);
   U4606 : NOR2X1 port map( A => n178, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b1);
   U4607 : NOR2X1 port map( A => n199, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b1);
   U4608 : NOR2X1 port map( A => n241, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b1);
   U4609 : NOR2X1 port map( A => n269, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b1);
   U4610 : NOR2X1 port map( A => n171, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b8);
   U4611 : NOR2X1 port map( A => n192, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b8);
   U4612 : NOR2X1 port map( A => n234, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b8);
   U4613 : NOR2X1 port map( A => n262, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b8);
   U4614 : NOR2X1 port map( A => n180, B => n173, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b6);
   U4615 : NOR2X1 port map( A => n201, B => n194, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b6);
   U4616 : NOR2X1 port map( A => n243, B => n236, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b6);
   U4617 : NOR2X1 port map( A => n271, B => n264, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b6);
   U4618 : NOR2X1 port map( A => n180, B => n172, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b7);
   U4619 : NOR2X1 port map( A => n201, B => n193, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b7);
   U4620 : NOR2X1 port map( A => n243, B => n235, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b7);
   U4621 : NOR2X1 port map( A => n271, B => n263, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b7);
   U4622 : NOR2X1 port map( A => n175, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b4);
   U4623 : NOR2X1 port map( A => n196, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b4);
   U4624 : NOR2X1 port map( A => n238, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b4);
   U4625 : NOR2X1 port map( A => n266, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b4);
   U4626 : NOR2X1 port map( A => n195, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b5);
   U4627 : NOR2X1 port map( A => n237, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b5);
   U4628 : NOR2X1 port map( A => n174, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b5);
   U4629 : NOR2X1 port map( A => n195, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b5);
   U4630 : NOR2X1 port map( A => n237, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b5);
   U4631 : NOR2X1 port map( A => n265, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b5);
   U4632 : NOR2X1 port map( A => n173, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b6);
   U4633 : NOR2X1 port map( A => n194, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b6);
   U4634 : NOR2X1 port map( A => n236, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b6);
   U4635 : NOR2X1 port map( A => n264, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b6);
   U4636 : NOR2X1 port map( A => n173, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b6);
   U4637 : NOR2X1 port map( A => n194, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b6);
   U4638 : NOR2X1 port map( A => n236, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b6);
   U4639 : NOR2X1 port map( A => n264, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b6);
   U4640 : NOR2X1 port map( A => n173, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b6);
   U4641 : NOR2X1 port map( A => n194, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b6);
   U4642 : NOR2X1 port map( A => n236, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b6);
   U4643 : NOR2X1 port map( A => n264, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b6);
   U4644 : NOR2X1 port map( A => n172, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b7);
   U4645 : NOR2X1 port map( A => n263, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b7);
   U4646 : NOR2X1 port map( A => n170, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b9);
   U4647 : NOR2X1 port map( A => n261, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b9);
   U4648 : NOR2X1 port map( A => n171, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b8);
   U4649 : NOR2X1 port map( A => n262, B => n278, Y => 
                           input_times_b0_mul_componentxUMxa2_and_b8);
   U4650 : NOR2X1 port map( A => n193, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b7);
   U4651 : NOR2X1 port map( A => n235, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b7);
   U4652 : NOR2X1 port map( A => n191, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b9);
   U4653 : NOR2X1 port map( A => n233, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b9);
   U4654 : NOR2X1 port map( A => n192, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b8);
   U4655 : NOR2X1 port map( A => n234, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b8);
   U4656 : NOR2X1 port map( A => n172, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b7);
   U4657 : NOR2X1 port map( A => n193, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b7);
   U4658 : NOR2X1 port map( A => n235, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b7);
   U4659 : NOR2X1 port map( A => n263, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b7);
   U4660 : NOR2X1 port map( A => n171, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b8);
   U4661 : NOR2X1 port map( A => n192, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b8);
   U4662 : NOR2X1 port map( A => n234, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b8);
   U4663 : NOR2X1 port map( A => n262, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b8);
   U4664 : NOR2X1 port map( A => n170, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b9);
   U4665 : NOR2X1 port map( A => n261, B => n275, Y => 
                           input_times_b0_mul_componentxUMxa5_and_b9);
   U4666 : NOR2X1 port map( A => n191, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b9);
   U4667 : NOR2X1 port map( A => n233, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b9);
   U4668 : NOR2X1 port map( A => n175, B => n4436, Y => 
                           input_p1_times_b1_mul_componentxUMxa13_and_b4);
   U4669 : NOR2X1 port map( A => n266, B => input_times_b0_mul_componentxn85, Y
                           => input_times_b0_mul_componentxUMxa13_and_b4);
   U4670 : NOR2X1 port map( A => n196, B => n4489, Y => 
                           input_p2_times_b2_mul_componentxUMxa13_and_b4);
   U4671 : NOR2X1 port map( A => n238, B => n4595, Y => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b4);
   U4672 : NOR2X1 port map( A => n179, B => n4433, Y => 
                           input_p1_times_b1_mul_componentxUMxa16_and_b0);
   U4673 : NOR2X1 port map( A => n270, B => input_times_b0_mul_componentxn82, Y
                           => input_times_b0_mul_componentxUMxa16_and_b0);
   U4674 : NOR2X1 port map( A => n200, B => n4486, Y => 
                           input_p2_times_b2_mul_componentxUMxa16_and_b0);
   U4675 : NOR2X1 port map( A => n242, B => n4592, Y => 
                           output_p2_times_a2_mul_componentxUMxa16_and_b0);
   U4676 : NOR2X1 port map( A => n179, B => n10, Y => 
                           input_p1_times_b1_mul_componentxUMxa17_and_b0);
   U4677 : XOR2X1 port map( A => n3687, B => input_previous_1_17_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_17_port);
   U4678 : NOR2X1 port map( A => n200, B => n11, Y => 
                           input_p2_times_b2_mul_componentxUMxa17_and_b0);
   U4679 : XOR2X1 port map( A => n3735, B => input_previous_2_17_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_17_port);
   U4680 : NOR2X1 port map( A => n242, B => n12, Y => 
                           output_p2_times_a2_mul_componentxUMxa17_and_b0);
   U4681 : XOR2X1 port map( A => n3831, B => output_previous_2_17_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_17_port);
   U4682 : NOR2X1 port map( A => n270, B => n13, Y => 
                           input_times_b0_mul_componentxUMxa17_and_b0);
   U4683 : XOR2X1 port map( A => n3639, B => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_17_port);
   U4684 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa15_and_b2,
                           B => input_p1_times_b1_mul_componentxUMxa16_and_b1, 
                           Y => n2718);
   U4685 : NOR2X1 port map( A => n177, B => n4434, Y => 
                           input_p1_times_b1_mul_componentxUMxa15_and_b2);
   U4686 : NOR2X1 port map( A => n178, B => n4433, Y => 
                           input_p1_times_b1_mul_componentxUMxa16_and_b1);
   U4687 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa14_and_b3,
                           B => n2717, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127715984_127849024_127850928);
   U4688 : NOR2X1 port map( A => n176, B => n4435, Y => 
                           input_p1_times_b1_mul_componentxUMxa14_and_b3);
   U4689 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa12_and_b5,
                           B => input_p1_times_b1_mul_componentxUMxa13_and_b4, 
                           Y => n2717);
   U4690 : NOR2X1 port map( A => n174, B => n4437, Y => 
                           input_p1_times_b1_mul_componentxUMxa12_and_b5);
   U4691 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa15_and_b2,
                           B => input_p2_times_b2_mul_componentxUMxa16_and_b1, 
                           Y => n2952);
   U4692 : NOR2X1 port map( A => n198, B => n4487, Y => 
                           input_p2_times_b2_mul_componentxUMxa15_and_b2);
   U4693 : NOR2X1 port map( A => n199, B => n4486, Y => 
                           input_p2_times_b2_mul_componentxUMxa16_and_b1);
   U4694 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa14_and_b3,
                           B => n2951, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127715984_127849024_127850928);
   U4695 : NOR2X1 port map( A => n197, B => n4488, Y => 
                           input_p2_times_b2_mul_componentxUMxa14_and_b3);
   U4696 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa12_and_b5,
                           B => input_p2_times_b2_mul_componentxUMxa13_and_b4, 
                           Y => n2951);
   U4697 : NOR2X1 port map( A => n195, B => n4490, Y => 
                           input_p2_times_b2_mul_componentxUMxa12_and_b5);
   U4698 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa15_and_b2
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa16_and_b1, Y =>
                           n3420);
   U4699 : NOR2X1 port map( A => n240, B => n4593, Y => 
                           output_p2_times_a2_mul_componentxUMxa15_and_b2);
   U4700 : NOR2X1 port map( A => n241, B => n4592, Y => 
                           output_p2_times_a2_mul_componentxUMxa16_and_b1);
   U4701 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa14_and_b3
                           , B => n3419, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127715984_127849024_127850928);
   U4702 : NOR2X1 port map( A => n239, B => n4594, Y => 
                           output_p2_times_a2_mul_componentxUMxa14_and_b3);
   U4703 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa12_and_b5
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa13_and_b4, Y =>
                           n3419);
   U4704 : NOR2X1 port map( A => n237, B => n4596, Y => 
                           output_p2_times_a2_mul_componentxUMxa12_and_b5);
   U4705 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa15_and_b2, B 
                           => input_times_b0_mul_componentxUMxa16_and_b1, Y => 
                           n2484);
   U4706 : NOR2X1 port map( A => n268, B => input_times_b0_mul_componentxn83, Y
                           => input_times_b0_mul_componentxUMxa15_and_b2);
   U4707 : NOR2X1 port map( A => n269, B => input_times_b0_mul_componentxn82, Y
                           => input_times_b0_mul_componentxUMxa16_and_b1);
   U4708 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa14_and_b3, B 
                           => n2483, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127715984_127849024_127850928);
   U4709 : NOR2X1 port map( A => n267, B => input_times_b0_mul_componentxn84, Y
                           => input_times_b0_mul_componentxUMxa14_and_b3);
   U4710 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa12_and_b5, B 
                           => input_times_b0_mul_componentxUMxa13_and_b4, Y => 
                           n2483);
   U4711 : NOR2X1 port map( A => n265, B => input_times_b0_mul_componentxn86, Y
                           => input_times_b0_mul_componentxUMxa12_and_b5);
   U4712 : NOR2X1 port map( A => n4421, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b11);
   U4713 : NOR2X1 port map( A => n4474, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b11);
   U4714 : NOR2X1 port map( A => n4580, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b11);
   U4715 : NOR2X1 port map( A => input_times_b0_mul_componentxn70, B => n276, Y
                           => input_times_b0_mul_componentxUMxa4_and_b11);
   U4716 : NOR2X1 port map( A => n4420, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b12);
   U4717 : NOR2X1 port map( A => n4473, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b12);
   U4718 : NOR2X1 port map( A => n4579, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b12);
   U4719 : NOR2X1 port map( A => input_times_b0_mul_componentxn69, B => n276, Y
                           => input_times_b0_mul_componentxUMxa4_and_b12);
   U4720 : NOR2X1 port map( A => input_times_b0_mul_componentxn68, B => n279, Y
                           => input_times_b0_mul_componentxUMxa1_and_b13);
   U4721 : NOR2X1 port map( A => n4419, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b13);
   U4722 : NOR2X1 port map( A => n4472, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b13);
   U4723 : NOR2X1 port map( A => n4578, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b13);
   U4724 : NOR2X1 port map( A => input_times_b0_mul_componentxn67, B => n279, Y
                           => input_times_b0_mul_componentxUMxa1_and_b14);
   U4725 : NOR2X1 port map( A => n4418, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b14);
   U4726 : NOR2X1 port map( A => n4471, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b14);
   U4727 : NOR2X1 port map( A => n4577, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b14);
   U4728 : NOR2X1 port map( A => n4417, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b15);
   U4729 : NOR2X1 port map( A => n4470, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b15);
   U4730 : NOR2X1 port map( A => n4576, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b15);
   U4731 : NOR2X1 port map( A => input_times_b0_mul_componentxn66, B => n279, Y
                           => input_times_b0_mul_componentxUMxa1_and_b15);
   U4732 : NOR2X1 port map( A => n192, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b8);
   U4733 : NOR2X1 port map( A => n234, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b8);
   U4734 : NOR2X1 port map( A => n170, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b9);
   U4735 : NOR2X1 port map( A => n191, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b9);
   U4736 : NOR2X1 port map( A => n233, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b9);
   U4737 : NOR2X1 port map( A => n261, B => n273, Y => 
                           input_times_b0_mul_componentxUMxa7_and_b9);
   U4738 : NOR2X1 port map( A => n4422, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b10);
   U4739 : NOR2X1 port map( A => n4475, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b10);
   U4740 : NOR2X1 port map( A => n4581, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b10);
   U4741 : NOR2X1 port map( A => input_times_b0_mul_componentxn71, B => n274, Y
                           => input_times_b0_mul_componentxUMxa6_and_b10);
   U4742 : NOR2X1 port map( A => n4422, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b10);
   U4743 : NOR2X1 port map( A => n4475, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b10);
   U4744 : NOR2X1 port map( A => n4581, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b10);
   U4745 : NOR2X1 port map( A => input_times_b0_mul_componentxn71, B => n275, Y
                           => input_times_b0_mul_componentxUMxa5_and_b10);
   U4746 : NOR2X1 port map( A => n4421, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b11);
   U4747 : NOR2X1 port map( A => n4474, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b11);
   U4748 : NOR2X1 port map( A => n4580, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b11);
   U4749 : NOR2X1 port map( A => input_times_b0_mul_componentxn70, B => n275, Y
                           => input_times_b0_mul_componentxUMxa5_and_b11);
   U4750 : NOR2X1 port map( A => n4420, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b12);
   U4751 : NOR2X1 port map( A => n4473, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b12);
   U4752 : NOR2X1 port map( A => n4579, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b12);
   U4753 : NOR2X1 port map( A => input_times_b0_mul_componentxn69, B => n277, Y
                           => input_times_b0_mul_componentxUMxa3_and_b12);
   U4754 : NOR2X1 port map( A => input_times_b0_mul_componentxn68, B => n277, Y
                           => input_times_b0_mul_componentxUMxa3_and_b13);
   U4755 : NOR2X1 port map( A => n4420, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b12);
   U4756 : NOR2X1 port map( A => n4473, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b12);
   U4757 : NOR2X1 port map( A => n4579, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b12);
   U4758 : NOR2X1 port map( A => input_times_b0_mul_componentxn69, B => n278, Y
                           => input_times_b0_mul_componentxUMxa2_and_b12);
   U4759 : NOR2X1 port map( A => n4419, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b13);
   U4760 : NOR2X1 port map( A => n4472, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b13);
   U4761 : NOR2X1 port map( A => n4578, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b13);
   U4762 : NOR2X1 port map( A => input_times_b0_mul_componentxn68, B => n278, Y
                           => input_times_b0_mul_componentxUMxa2_and_b13);
   U4763 : NOR2X1 port map( A => n4419, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b13);
   U4764 : NOR2X1 port map( A => n4472, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b13);
   U4765 : NOR2X1 port map( A => n4578, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b13);
   U4766 : NOR2X1 port map( A => n280, B => input_times_b0_mul_componentxn67, Y
                           => input_times_b0_mul_componentxUMxa0_and_b14);
   U4767 : NOR2X1 port map( A => n189, B => n4418, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b14);
   U4768 : NOR2X1 port map( A => n210, B => n4471, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b14);
   U4769 : NOR2X1 port map( A => n252, B => n4577, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b14);
   U4770 : NOR2X1 port map( A => n189, B => n4417, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b15);
   U4771 : NOR2X1 port map( A => n210, B => n4470, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b15);
   U4772 : NOR2X1 port map( A => n252, B => n4576, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b15);
   U4773 : NOR2X1 port map( A => n280, B => input_times_b0_mul_componentxn66, Y
                           => input_times_b0_mul_componentxUMxa0_and_b15);
   U4774 : NOR2X1 port map( A => n189, B => n4416, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b16);
   U4775 : NOR2X1 port map( A => n210, B => n4469, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b16);
   U4776 : NOR2X1 port map( A => n252, B => n4575, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b16);
   U4777 : NOR2X1 port map( A => n280, B => input_times_b0_mul_componentxn65, Y
                           => input_times_b0_mul_componentxUMxa0_and_b16);
   U4778 : NOR2X1 port map( A => n170, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b9);
   U4779 : NOR2X1 port map( A => n261, B => n274, Y => 
                           input_times_b0_mul_componentxUMxa6_and_b9);
   U4780 : NOR2X1 port map( A => n191, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b9);
   U4781 : NOR2X1 port map( A => n233, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b9);
   U4782 : NOR2X1 port map( A => n172, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b7);
   U4783 : NOR2X1 port map( A => n193, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b7);
   U4784 : NOR2X1 port map( A => n235, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b7);
   U4785 : NOR2X1 port map( A => n263, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b7);
   U4786 : NOR2X1 port map( A => n171, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b8);
   U4787 : NOR2X1 port map( A => n192, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b8);
   U4788 : NOR2X1 port map( A => n234, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b8);
   U4789 : NOR2X1 port map( A => n262, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b8);
   U4790 : NOR2X1 port map( A => n189, B => n178, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b1);
   U4791 : NOR2X1 port map( A => n280, B => n269, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b1);
   U4792 : NOR2X1 port map( A => n210, B => n199, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b1);
   U4793 : NOR2X1 port map( A => n252, B => n241, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b1);
   U4794 : NOR2X1 port map( A => n179, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b0);
   U4795 : NOR2X1 port map( A => n200, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b0);
   U4796 : NOR2X1 port map( A => n242, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b0);
   U4797 : NOR2X1 port map( A => n270, B => n279, Y => 
                           input_times_b0_mul_componentxUMxa1_and_b0);
   U4798 : NOR2X1 port map( A => n173, B => n4438, Y => 
                           input_p1_times_b1_mul_componentxUMxa11_and_b6);
   U4799 : NOR2X1 port map( A => n264, B => input_times_b0_mul_componentxn87, Y
                           => input_times_b0_mul_componentxUMxa11_and_b6);
   U4800 : NOR2X1 port map( A => n194, B => n4491, Y => 
                           input_p2_times_b2_mul_componentxUMxa11_and_b6);
   U4801 : NOR2X1 port map( A => n236, B => n4597, Y => 
                           output_p2_times_a2_mul_componentxUMxa11_and_b6);
   U4802 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa9_and_b8, 
                           B => input_p1_times_b1_mul_componentxUMxa10_and_b7, 
                           Y => n2716);
   U4803 : NOR2X1 port map( A => n180, B => n171, Y => 
                           input_p1_times_b1_mul_componentxUMxa9_and_b8);
   U4804 : NOR2X1 port map( A => n172, B => n4439, Y => 
                           input_p1_times_b1_mul_componentxUMxa10_and_b7);
   U4805 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa9_and_b8, 
                           B => input_p2_times_b2_mul_componentxUMxa10_and_b7, 
                           Y => n2950);
   U4806 : NOR2X1 port map( A => n201, B => n192, Y => 
                           input_p2_times_b2_mul_componentxUMxa9_and_b8);
   U4807 : NOR2X1 port map( A => n193, B => n4492, Y => 
                           input_p2_times_b2_mul_componentxUMxa10_and_b7);
   U4808 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa9_and_b8,
                           B => output_p2_times_a2_mul_componentxUMxa10_and_b7,
                           Y => n3418);
   U4809 : NOR2X1 port map( A => n243, B => n234, Y => 
                           output_p2_times_a2_mul_componentxUMxa9_and_b8);
   U4810 : NOR2X1 port map( A => n235, B => n4598, Y => 
                           output_p2_times_a2_mul_componentxUMxa10_and_b7);
   U4811 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa9_and_b8, B 
                           => input_times_b0_mul_componentxUMxa10_and_b7, Y => 
                           n2482);
   U4812 : NOR2X1 port map( A => n271, B => n262, Y => 
                           input_times_b0_mul_componentxUMxa9_and_b8);
   U4813 : NOR2X1 port map( A => n263, B => input_times_b0_mul_componentxn88, Y
                           => input_times_b0_mul_componentxUMxa10_and_b7);
   U4814 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa6_and_b11,
                           B => input_p1_times_b1_mul_componentxUMxa7_and_b10, 
                           Y => n2715);
   U4815 : NOR2X1 port map( A => n4421, B => n183, Y => 
                           input_p1_times_b1_mul_componentxUMxa6_and_b11);
   U4816 : NOR2X1 port map( A => n4422, B => n182, Y => 
                           input_p1_times_b1_mul_componentxUMxa7_and_b10);
   U4817 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa6_and_b11,
                           B => input_p2_times_b2_mul_componentxUMxa7_and_b10, 
                           Y => n2949);
   U4818 : NOR2X1 port map( A => n4474, B => n204, Y => 
                           input_p2_times_b2_mul_componentxUMxa6_and_b11);
   U4819 : NOR2X1 port map( A => n4475, B => n203, Y => 
                           input_p2_times_b2_mul_componentxUMxa7_and_b10);
   U4820 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa6_and_b11
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b10, Y =>
                           n3417);
   U4821 : NOR2X1 port map( A => n4580, B => n246, Y => 
                           output_p2_times_a2_mul_componentxUMxa6_and_b11);
   U4822 : NOR2X1 port map( A => n4581, B => n245, Y => 
                           output_p2_times_a2_mul_componentxUMxa7_and_b10);
   U4823 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa6_and_b11, B 
                           => input_times_b0_mul_componentxUMxa7_and_b10, Y => 
                           n2481);
   U4824 : NOR2X1 port map( A => input_times_b0_mul_componentxn70, B => n274, Y
                           => input_times_b0_mul_componentxUMxa6_and_b11);
   U4825 : NOR2X1 port map( A => input_times_b0_mul_componentxn71, B => n273, Y
                           => input_times_b0_mul_componentxUMxa7_and_b10);
   U4826 : NOR2X1 port map( A => n189, B => n179, Y => 
                           input_p1_times_b1_mul_componentxUMxfirst_vector_0_port);
   U4827 : NOR2X1 port map( A => n210, B => n200, Y => 
                           input_p2_times_b2_mul_componentxUMxfirst_vector_0_port);
   U4828 : NOR2X1 port map( A => n252, B => n242, Y => 
                           output_p2_times_a2_mul_componentxUMxfirst_vector_0_port);
   U4829 : NOR2X1 port map( A => n280, B => n270, Y => 
                           input_times_b0_mul_componentxUMxfirst_vector_0_port)
                           ;
   U4830 : NOR2X1 port map( A => input_times_b0_mul_componentxn67, B => n278, Y
                           => input_times_b0_mul_componentxUMxa2_and_b14);
   U4831 : NOR2X1 port map( A => n4418, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b14);
   U4832 : NOR2X1 port map( A => n4471, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b14);
   U4833 : NOR2X1 port map( A => n4577, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b14);
   U4834 : NOR2X1 port map( A => input_times_b0_mul_componentxn68, B => n276, Y
                           => input_times_b0_mul_componentxUMxa4_and_b13);
   U4835 : NOR2X1 port map( A => n4419, B => n185, Y => 
                           input_p1_times_b1_mul_componentxUMxa4_and_b13);
   U4836 : NOR2X1 port map( A => n4472, B => n206, Y => 
                           input_p2_times_b2_mul_componentxUMxa4_and_b13);
   U4837 : NOR2X1 port map( A => n4578, B => n248, Y => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b13);
   U4838 : NOR2X1 port map( A => n4417, B => n187, Y => 
                           input_p1_times_b1_mul_componentxUMxa2_and_b15);
   U4839 : NOR2X1 port map( A => n4470, B => n208, Y => 
                           input_p2_times_b2_mul_componentxUMxa2_and_b15);
   U4840 : NOR2X1 port map( A => n4576, B => n250, Y => 
                           output_p2_times_a2_mul_componentxUMxa2_and_b15);
   U4841 : NOR2X1 port map( A => input_times_b0_mul_componentxn66, B => n278, Y
                           => input_times_b0_mul_componentxUMxa2_and_b15);
   U4842 : NOR2X1 port map( A => n170, B => n181, Y => 
                           input_p1_times_b1_mul_componentxUMxa8_and_b9);
   U4843 : NOR2X1 port map( A => n191, B => n202, Y => 
                           input_p2_times_b2_mul_componentxUMxa8_and_b9);
   U4844 : NOR2X1 port map( A => n233, B => n244, Y => 
                           output_p2_times_a2_mul_componentxUMxa8_and_b9);
   U4845 : NOR2X1 port map( A => n261, B => n272, Y => 
                           input_times_b0_mul_componentxUMxa8_and_b9);
   U4846 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa0_and_b17,
                           B => input_p1_times_b1_mul_componentxUMxa1_and_b16, 
                           Y => n2713);
   U4847 : NOR2X1 port map( A => n189, B => n21, Y => 
                           input_p1_times_b1_mul_componentxUMxa0_and_b17);
   U4848 : NOR2X1 port map( A => n4416, B => n188, Y => 
                           input_p1_times_b1_mul_componentxUMxa1_and_b16);
   U4849 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa0_and_b17,
                           B => input_p2_times_b2_mul_componentxUMxa1_and_b16, 
                           Y => n2947);
   U4850 : NOR2X1 port map( A => n210, B => n22, Y => 
                           input_p2_times_b2_mul_componentxUMxa0_and_b17);
   U4851 : NOR2X1 port map( A => n4469, B => n209, Y => 
                           input_p2_times_b2_mul_componentxUMxa1_and_b16);
   U4852 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa0_and_b17
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b16, Y =>
                           n3415);
   U4853 : NOR2X1 port map( A => n252, B => n23, Y => 
                           output_p2_times_a2_mul_componentxUMxa0_and_b17);
   U4854 : NOR2X1 port map( A => n4575, B => n251, Y => 
                           output_p2_times_a2_mul_componentxUMxa1_and_b16);
   U4855 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa0_and_b17, B 
                           => input_times_b0_mul_componentxUMxa1_and_b16, Y => 
                           n2479);
   U4856 : NOR2X1 port map( A => n280, B => n24, Y => 
                           input_times_b0_mul_componentxUMxa0_and_b17);
   U4857 : NOR2X1 port map( A => input_times_b0_mul_componentxn65, B => n279, Y
                           => input_times_b0_mul_componentxUMxa1_and_b16);
   U4858 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa5_and_b12,
                           B => n2714, Y => 
                           input_p1_times_b1_mul_componentxUMxsum_layer1_127674016_127675920_127731136);
   U4859 : NOR2X1 port map( A => n4420, B => n184, Y => 
                           input_p1_times_b1_mul_componentxUMxa5_and_b12);
   U4860 : XOR2X1 port map( A => input_p1_times_b1_mul_componentxUMxa3_and_b14,
                           B => input_p1_times_b1_mul_componentxUMxa4_and_b13, 
                           Y => n2714);
   U4861 : NOR2X1 port map( A => n4418, B => n186, Y => 
                           input_p1_times_b1_mul_componentxUMxa3_and_b14);
   U4862 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa5_and_b12,
                           B => n2948, Y => 
                           input_p2_times_b2_mul_componentxUMxsum_layer1_127674016_127675920_127731136);
   U4863 : NOR2X1 port map( A => n4473, B => n205, Y => 
                           input_p2_times_b2_mul_componentxUMxa5_and_b12);
   U4864 : XOR2X1 port map( A => input_p2_times_b2_mul_componentxUMxa3_and_b14,
                           B => input_p2_times_b2_mul_componentxUMxa4_and_b13, 
                           Y => n2948);
   U4865 : NOR2X1 port map( A => n4471, B => n207, Y => 
                           input_p2_times_b2_mul_componentxUMxa3_and_b14);
   U4866 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa5_and_b12
                           , B => n3416, Y => 
                           output_p2_times_a2_mul_componentxUMxsum_layer1_127674016_127675920_127731136);
   U4867 : NOR2X1 port map( A => n4579, B => n247, Y => 
                           output_p2_times_a2_mul_componentxUMxa5_and_b12);
   U4868 : XOR2X1 port map( A => output_p2_times_a2_mul_componentxUMxa3_and_b14
                           , B => 
                           output_p2_times_a2_mul_componentxUMxa4_and_b13, Y =>
                           n3416);
   U4869 : NOR2X1 port map( A => n4577, B => n249, Y => 
                           output_p2_times_a2_mul_componentxUMxa3_and_b14);
   U4870 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa5_and_b12, B 
                           => n2480, Y => 
                           input_times_b0_mul_componentxUMxsum_layer1_127674016_127675920_127731136);
   U4871 : NOR2X1 port map( A => input_times_b0_mul_componentxn69, B => n275, Y
                           => input_times_b0_mul_componentxUMxa5_and_b12);
   U4872 : XOR2X1 port map( A => input_times_b0_mul_componentxUMxa3_and_b14, B 
                           => input_times_b0_mul_componentxUMxa4_and_b13, Y => 
                           n2480);
   U4873 : NOR2X1 port map( A => input_times_b0_mul_componentxn67, B => n277, Y
                           => input_times_b0_mul_componentxUMxa3_and_b14);
   U4874 : OAI2BB2X1 port map( B0 => n1174, B1 => n319, A0N => 
                           input_previous_0_17_port, A1N => n320, Y => 
                           input_prev_0_registerxn20);
   U4875 : OR2X2 port map( A => n367, B => change_input_port, Y => n103);
   U4876 : INVX1 port map( A => n103, Y => n1870);
   U4877 : OR2X2 port map( A => n367, B => change_input_port, Y => n104);
   U4878 : INVX1 port map( A => n104, Y => n1980);
   U4879 : OR2X2 port map( A => n368, B => change_input_port, Y => n105);
   U4880 : INVX1 port map( A => n105, Y => n2089);
   U4881 : OR2X2 port map( A => n368, B => change_input_port, Y => n106);
   U4882 : INVX1 port map( A => n106, Y => n2199);
   U4883 : OR2X2 port map( A => n367, B => change_input_port, Y => n107);
   U4884 : INVX1 port map( A => n107, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn3);
   U4885 : INVX1 port map( A => change_input_port, Y => n1260);
   U4886 : INVX1 port map( A => n4203, Y => n374);
   U4887 : INVX1 port map( A => n4259, Y => n376);
   U4888 : INVX1 port map( A => n4369, Y => n378);
   U4889 : INVX1 port map( A => input_times_b0_div_componentxn24, Y => n380);
   U4890 : AOI22X1 port map( A0 => n335, A1 => n338, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_10_port, 
                           B1 => n336, Y => n4422);
   U4891 : XOR2X1 port map( A => n3710, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_10_port);
   U4892 : NAND2X1 port map( A => n3695, B => n337, Y => n3710);
   U4893 : AOI22X1 port map( A0 => n326, A1 => n329, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_10_port, 
                           B1 => n327, Y => n4475);
   U4894 : XOR2X1 port map( A => n3758, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_10_port);
   U4895 : NAND2X1 port map( A => n3743, B => n328, Y => n3758);
   U4896 : AOI22X1 port map( A0 => n362, A1 => n365, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_10_port, 
                           B1 => n363, Y => n4528);
   U4897 : XOR2X1 port map( A => n3806, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_10_port);
   U4898 : NAND2X1 port map( A => n3791, B => n364, Y => n3806);
   U4899 : AOI22X1 port map( A0 => n353, A1 => n356, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_10_port, 
                           B1 => n354, Y => n4581);
   U4900 : XOR2X1 port map( A => n3854, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_10_port);
   U4901 : NAND2X1 port map( A => n3839, B => n355, Y => n3854);
   U4902 : AOI22X1 port map( A0 => n344, A1 => n347, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_10_port, 
                           B1 => n345, Y => input_times_b0_mul_componentxn71);
   U4903 : XOR2X1 port map( A => n3662, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_10_port);
   U4904 : NAND2X1 port map( A => n3647, B => n346, Y => n3662);
   U4905 : AOI22X1 port map( A0 => n362, A1 => n365, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_11_port, 
                           B1 => n363, Y => n4527);
   U4906 : XOR2X1 port map( A => n3804, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_11_port);
   U4907 : AOI22X1 port map( A0 => n335, A1 => n338, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_11_port, 
                           B1 => n336, Y => n4421);
   U4908 : XOR2X1 port map( A => n3708, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_11_port);
   U4909 : AOI22X1 port map( A0 => n326, A1 => n329, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_11_port, 
                           B1 => n327, Y => n4474);
   U4910 : XOR2X1 port map( A => n3756, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_11_port);
   U4911 : AOI22X1 port map( A0 => n353, A1 => n356, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_11_port, 
                           B1 => n354, Y => n4580);
   U4912 : XOR2X1 port map( A => n3852, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_11_port);
   U4913 : AOI22X1 port map( A0 => n344, A1 => n347, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_11_port, 
                           B1 => n345, Y => input_times_b0_mul_componentxn70);
   U4914 : XOR2X1 port map( A => n3660, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_11_port);
   U4915 : AOI22X1 port map( A0 => n362, A1 => n364, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_12_port, 
                           B1 => n363, Y => n4526);
   U4916 : XOR2X1 port map( A => n3805, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_12_port);
   U4917 : OR2X2 port map( A => n3804, B => n363, Y => n3805);
   U4918 : AOI22X1 port map( A0 => n335, A1 => n338, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_12_port, 
                           B1 => n336, Y => n4420);
   U4919 : XOR2X1 port map( A => n3709, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_12_port);
   U4920 : OR2X2 port map( A => n3708, B => n336, Y => n3709);
   U4921 : AOI22X1 port map( A0 => n326, A1 => n329, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_12_port, 
                           B1 => n327, Y => n4473);
   U4922 : XOR2X1 port map( A => n3757, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_12_port);
   U4923 : OR2X2 port map( A => n3756, B => n327, Y => n3757);
   U4924 : AOI22X1 port map( A0 => n353, A1 => n356, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_12_port, 
                           B1 => n354, Y => n4579);
   U4925 : XOR2X1 port map( A => n3853, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_12_port);
   U4926 : OR2X2 port map( A => n3852, B => n354, Y => n3853);
   U4927 : AOI22X1 port map( A0 => n344, A1 => n347, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_12_port, 
                           B1 => n345, Y => input_times_b0_mul_componentxn69);
   U4928 : XOR2X1 port map( A => n3661, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_12_port);
   U4929 : OR2X2 port map( A => n3660, B => n345, Y => n3661);
   U4930 : AOI22X1 port map( A0 => n341, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_9_port
                           , B1 => parameter_B0_div(7), Y => 
                           input_times_b0_div_componentxn54);
   U4931 : XNOR2X1 port map( A => n3882, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_9_port
                           );
   U4932 : AOI22X1 port map( A0 => n332, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_9_port, 
                           B1 => parameter_B1_div(7), Y => n4232);
   U4933 : XNOR2X1 port map( A => n3925, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_9_port);
   U4934 : AOI22X1 port map( A0 => n323, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_9_port, 
                           B1 => parameter_B2_div(7), Y => n4288);
   U4935 : XNOR2X1 port map( A => n3968, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_9_port);
   U4936 : AOI22X1 port map( A0 => n359, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_9_port, 
                           B1 => parameter_A1_div(7), Y => n4342);
   U4937 : XNOR2X1 port map( A => n4011, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_9_port);
   U4938 : AOI22X1 port map( A0 => n350, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_9_port, 
                           B1 => parameter_A2_div(7), Y => n4398);
   U4939 : XNOR2X1 port map( A => n4054, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_9_port);
   U4940 : AOI22X1 port map( A0 => n343, A1 => n348, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_13_port, 
                           B1 => n344, Y => input_times_b0_mul_componentxn68);
   U4941 : XOR2X1 port map( A => n3658, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_13_port);
   U4942 : AOI22X1 port map( A0 => n335, A1 => n339, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_13_port, 
                           B1 => n336, Y => n4419);
   U4943 : XOR2X1 port map( A => n3706, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_13_port);
   U4944 : AOI22X1 port map( A0 => n326, A1 => n330, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_13_port, 
                           B1 => n327, Y => n4472);
   U4945 : XOR2X1 port map( A => n3754, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_13_port);
   U4946 : AOI22X1 port map( A0 => n362, A1 => n364, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_13_port, 
                           B1 => n363, Y => n4525);
   U4947 : XOR2X1 port map( A => n3802, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_13_port);
   U4948 : AOI22X1 port map( A0 => n353, A1 => n357, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_13_port, 
                           B1 => n354, Y => n4578);
   U4949 : XOR2X1 port map( A => n3850, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_13_port);
   U4950 : AOI22X1 port map( A0 => n344, A1 => n348, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_14_port, 
                           B1 => n344, Y => input_times_b0_mul_componentxn67);
   U4951 : XOR2X1 port map( A => n3659, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_14_port);
   U4952 : OR2X2 port map( A => n345, B => n3658, Y => n3659);
   U4953 : AOI22X1 port map( A0 => n335, A1 => n339, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_14_port, 
                           B1 => n336, Y => n4418);
   U4954 : XOR2X1 port map( A => n3707, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_14_port);
   U4955 : OR2X2 port map( A => n336, B => n3706, Y => n3707);
   U4956 : AOI22X1 port map( A0 => n326, A1 => n330, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_14_port, 
                           B1 => n327, Y => n4471);
   U4957 : XOR2X1 port map( A => n3755, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_14_port);
   U4958 : OR2X2 port map( A => n327, B => n3754, Y => n3755);
   U4959 : AOI22X1 port map( A0 => n362, A1 => n366, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_14_port, 
                           B1 => n363, Y => n4524);
   U4960 : XOR2X1 port map( A => n3803, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_14_port);
   U4961 : OR2X2 port map( A => n363, B => n3802, Y => n3803);
   U4962 : AOI22X1 port map( A0 => n353, A1 => n357, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_14_port, 
                           B1 => n354, Y => n4577);
   U4963 : XOR2X1 port map( A => n3851, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_14_port);
   U4964 : OR2X2 port map( A => n354, B => n3850, Y => n3851);
   U4965 : AOI22X1 port map( A0 => n335, A1 => n337, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_15_port, 
                           B1 => n335, Y => n4417);
   U4966 : XNOR2X1 port map( A => n3705, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_15_port);
   U4967 : AOI22X1 port map( A0 => n326, A1 => n328, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_15_port, 
                           B1 => n326, Y => n4470);
   U4968 : XNOR2X1 port map( A => n3753, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_15_port);
   U4969 : AOI22X1 port map( A0 => n362, A1 => n364, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_15_port, 
                           B1 => n362, Y => n4523);
   U4970 : XNOR2X1 port map( A => n3801, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_15_port);
   U4971 : AOI22X1 port map( A0 => n353, A1 => n355, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_15_port, 
                           B1 => n353, Y => n4576);
   U4972 : XNOR2X1 port map( A => n3849, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_15_port);
   U4973 : AOI22X1 port map( A0 => n343, A1 => n346, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_15_port, 
                           B1 => n345, Y => input_times_b0_mul_componentxn66);
   U4974 : XNOR2X1 port map( A => n3657, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_15_port);
   U4975 : AOI22X1 port map( A0 => n341, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_8_port
                           , B1 => n341, Y => input_times_b0_div_componentxn53)
                           ;
   U4976 : XOR2X1 port map( A => n3883, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_8_port
                           );
   U4977 : OR2X2 port map( A => parameter_B0_div(7), B => n3884, Y => n3883);
   U4978 : AOI22X1 port map( A0 => n332, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_8_port, 
                           B1 => n332, Y => n4231);
   U4979 : XOR2X1 port map( A => n3926, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_8_port);
   U4980 : OR2X2 port map( A => parameter_B1_div(7), B => n3927, Y => n3926);
   U4981 : AOI22X1 port map( A0 => n323, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_8_port, 
                           B1 => n323, Y => n4287);
   U4982 : XOR2X1 port map( A => n3969, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_8_port);
   U4983 : OR2X2 port map( A => parameter_B2_div(7), B => n3970, Y => n3969);
   U4984 : AOI22X1 port map( A0 => n359, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_8_port, 
                           B1 => n359, Y => n4341);
   U4985 : XOR2X1 port map( A => n4012, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_8_port);
   U4986 : OR2X2 port map( A => parameter_A1_div(7), B => n4013, Y => n4012);
   U4987 : AOI22X1 port map( A0 => n350, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_8_port, 
                           B1 => n350, Y => n4397);
   U4988 : XOR2X1 port map( A => n4055, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_8_port);
   U4989 : OR2X2 port map( A => parameter_A2_div(7), B => n4056, Y => n4055);
   U4990 : AOI22X1 port map( A0 => n362, A1 => n364, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_16_port, 
                           B1 => n362, Y => n4522);
   U4991 : XNOR2X1 port map( A => n3800, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_16_port);
   U4992 : AOI22X1 port map( A0 => n335, A1 => n337, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_16_port, 
                           B1 => n335, Y => n4416);
   U4993 : XNOR2X1 port map( A => n3704, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_16_port);
   U4994 : AOI22X1 port map( A0 => n326, A1 => n328, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_16_port, 
                           B1 => n326, Y => n4469);
   U4995 : XNOR2X1 port map( A => n3752, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_16_port);
   U4996 : AOI22X1 port map( A0 => n353, A1 => n355, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_16_port, 
                           B1 => n353, Y => n4575);
   U4997 : XNOR2X1 port map( A => n3848, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_16_port);
   U4998 : AOI22X1 port map( A0 => n344, A1 => n346, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_16_port, 
                           B1 => n344, Y => input_times_b0_mul_componentxn65);
   U4999 : XNOR2X1 port map( A => n3656, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_16_port);
   U5000 : AOI22X1 port map( A0 => n341, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_7_port
                           , B1 => n341, Y => input_times_b0_div_componentxn52)
                           ;
   U5001 : XOR2X1 port map( A => n3884, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_7_port
                           );
   U5002 : AOI22X1 port map( A0 => n332, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_7_port, 
                           B1 => n332, Y => n4230);
   U5003 : XOR2X1 port map( A => n3927, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_7_port);
   U5004 : AOI22X1 port map( A0 => n323, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_7_port, 
                           B1 => n323, Y => n4286);
   U5005 : XOR2X1 port map( A => n3970, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_7_port);
   U5006 : AOI22X1 port map( A0 => n359, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_7_port, 
                           B1 => n359, Y => n4340);
   U5007 : XOR2X1 port map( A => n4013, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_7_port);
   U5008 : AOI22X1 port map( A0 => n350, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_7_port, 
                           B1 => n350, Y => n4396);
   U5009 : XOR2X1 port map( A => n4056, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_7_port);
   U5010 : AOI22X1 port map( A0 => n341, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_11_port, 
                           B1 => n341, Y => input_times_b0_div_componentxn56);
   U5011 : XOR2X1 port map( A => n3895, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_11_port);
   U5012 : AOI22X1 port map( A0 => n332, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_11_port, 
                           B1 => n332, Y => n4234);
   U5013 : XOR2X1 port map( A => n3938, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_11_port);
   U5014 : AOI22X1 port map( A0 => n323, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_11_port, 
                           B1 => n323, Y => n4290);
   U5015 : XOR2X1 port map( A => n3981, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_11_port);
   U5016 : AOI22X1 port map( A0 => n359, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_11_port, 
                           B1 => n359, Y => n4344);
   U5017 : XOR2X1 port map( A => n4024, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_11_port);
   U5018 : AOI22X1 port map( A0 => n350, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_11_port, 
                           B1 => n350, Y => n4400);
   U5019 : XOR2X1 port map( A => n4067, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_11_port);
   U5020 : AOI22X1 port map( A0 => n341, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_13_port, 
                           B1 => n341, Y => input_times_b0_div_componentxn58);
   U5021 : XOR2X1 port map( A => n3893, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_13_port);
   U5022 : AOI22X1 port map( A0 => n332, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_13_port, 
                           B1 => n332, Y => n4236);
   U5023 : XOR2X1 port map( A => n3936, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_13_port);
   U5024 : AOI22X1 port map( A0 => n323, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_13_port, 
                           B1 => n323, Y => n4292);
   U5025 : XOR2X1 port map( A => n3979, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_13_port);
   U5026 : AOI22X1 port map( A0 => n359, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_13_port, 
                           B1 => n359, Y => n4346);
   U5027 : XOR2X1 port map( A => n4022, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_13_port);
   U5028 : AOI22X1 port map( A0 => n350, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_13_port, 
                           B1 => n350, Y => n4402);
   U5029 : XOR2X1 port map( A => n4065, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_13_port);
   U5030 : AOI22X1 port map( A0 => n341, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_10_port, 
                           B1 => parameter_B0_div(7), Y => 
                           input_times_b0_div_componentxn55);
   U5031 : XOR2X1 port map( A => n3897, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_10_port);
   U5032 : NAND2X1 port map( A => n3882, B => n342, Y => n3897);
   U5033 : AOI22X1 port map( A0 => n332, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_10_port, 
                           B1 => parameter_B1_div(7), Y => n4233);
   U5034 : XOR2X1 port map( A => n3940, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_10_port);
   U5035 : NAND2X1 port map( A => n3925, B => n333, Y => n3940);
   U5036 : AOI22X1 port map( A0 => n323, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_10_port, 
                           B1 => parameter_B2_div(7), Y => n4289);
   U5037 : XOR2X1 port map( A => n3983, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_10_port);
   U5038 : NAND2X1 port map( A => n3968, B => n324, Y => n3983);
   U5039 : AOI22X1 port map( A0 => n359, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_10_port, 
                           B1 => parameter_A1_div(7), Y => n4343);
   U5040 : XOR2X1 port map( A => n4026, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_10_port);
   U5041 : NAND2X1 port map( A => n4011, B => n360, Y => n4026);
   U5042 : AOI22X1 port map( A0 => n350, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_10_port, 
                           B1 => parameter_A2_div(7), Y => n4399);
   U5043 : XOR2X1 port map( A => n4069, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_10_port);
   U5044 : NAND2X1 port map( A => n4054, B => n351, Y => n4069);
   U5045 : AOI22X1 port map( A0 => n341, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_12_port, 
                           B1 => parameter_B0_div(7), Y => 
                           input_times_b0_div_componentxn57);
   U5046 : XOR2X1 port map( A => n3896, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_12_port);
   U5047 : OR2X2 port map( A => n3895, B => parameter_B0_div(7), Y => n3896);
   U5048 : AOI22X1 port map( A0 => n332, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_12_port, 
                           B1 => parameter_B1_div(7), Y => n4235);
   U5049 : XOR2X1 port map( A => n3939, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_12_port);
   U5050 : OR2X2 port map( A => n3938, B => parameter_B1_div(7), Y => n3939);
   U5051 : AOI22X1 port map( A0 => n323, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_12_port, 
                           B1 => parameter_B2_div(7), Y => n4291);
   U5052 : XOR2X1 port map( A => n3982, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_12_port);
   U5053 : OR2X2 port map( A => n3981, B => parameter_B2_div(7), Y => n3982);
   U5054 : AOI22X1 port map( A0 => n359, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_12_port, 
                           B1 => parameter_A1_div(7), Y => n4345);
   U5055 : XOR2X1 port map( A => n4025, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_12_port);
   U5056 : OR2X2 port map( A => n4024, B => parameter_A1_div(7), Y => n4025);
   U5057 : AOI22X1 port map( A0 => n350, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_12_port, 
                           B1 => parameter_A2_div(7), Y => n4401);
   U5058 : XOR2X1 port map( A => n4068, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_12_port);
   U5059 : OR2X2 port map( A => n4067, B => parameter_A2_div(7), Y => n4068);
   U5060 : AOI22X1 port map( A0 => n340, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_14_port, 
                           B1 => parameter_B0_div(7), Y => 
                           input_times_b0_div_componentxn59);
   U5061 : XOR2X1 port map( A => n3894, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_14_port);
   U5062 : OR2X2 port map( A => parameter_B0_div(7), B => n3893, Y => n3894);
   U5063 : AOI22X1 port map( A0 => n331, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_14_port, 
                           B1 => parameter_B1_div(7), Y => n4237);
   U5064 : XOR2X1 port map( A => n3937, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_14_port);
   U5065 : OR2X2 port map( A => parameter_B1_div(7), B => n3936, Y => n3937);
   U5066 : AOI22X1 port map( A0 => n322, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_14_port, 
                           B1 => parameter_B2_div(7), Y => n4293);
   U5067 : XOR2X1 port map( A => n3980, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_14_port);
   U5068 : OR2X2 port map( A => parameter_B2_div(7), B => n3979, Y => n3980);
   U5069 : AOI22X1 port map( A0 => n358, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_14_port, 
                           B1 => parameter_A1_div(7), Y => n4347);
   U5070 : XOR2X1 port map( A => n4023, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_14_port);
   U5071 : OR2X2 port map( A => parameter_A1_div(7), B => n4022, Y => n4023);
   U5072 : AOI22X1 port map( A0 => n349, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_14_port, 
                           B1 => parameter_A2_div(7), Y => n4403);
   U5073 : XOR2X1 port map( A => n4066, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_14_port);
   U5074 : OR2X2 port map( A => parameter_A2_div(7), B => n4065, Y => n4066);
   U5075 : AOI22X1 port map( A0 => n340, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_15_port, 
                           B1 => parameter_B0_div(7), Y => 
                           input_times_b0_div_componentxn60);
   U5076 : XNOR2X1 port map( A => n3892, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_15_port);
   U5077 : AOI22X1 port map( A0 => n331, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_15_port, 
                           B1 => parameter_B1_div(7), Y => n4238);
   U5078 : XNOR2X1 port map( A => n3935, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_15_port);
   U5079 : AOI22X1 port map( A0 => n322, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_15_port, 
                           B1 => parameter_B2_div(7), Y => n4294);
   U5080 : XNOR2X1 port map( A => n3978, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_15_port);
   U5081 : AOI22X1 port map( A0 => n358, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_15_port, 
                           B1 => parameter_A1_div(7), Y => n4348);
   U5082 : XNOR2X1 port map( A => n4021, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_15_port);
   U5083 : AOI22X1 port map( A0 => n349, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_15_port, 
                           B1 => parameter_A2_div(7), Y => n4404);
   U5084 : XNOR2X1 port map( A => n4064, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_15_port);
   U5085 : NOR2X1 port map( A => n336, B => n3697, Y => n3695);
   U5086 : NOR2X1 port map( A => n327, B => n3745, Y => n3743);
   U5087 : NOR2X1 port map( A => n363, B => n3793, Y => n3791);
   U5088 : NOR2X1 port map( A => n354, B => n3841, Y => n3839);
   U5089 : NOR2X1 port map( A => n345, B => n3649, Y => n3647);
   U5090 : NOR2X1 port map( A => parameter_B0_div(7), B => n3884, Y => n3882);
   U5091 : NOR2X1 port map( A => parameter_B1_div(7), B => n3927, Y => n3925);
   U5092 : NOR2X1 port map( A => parameter_B2_div(7), B => n3970, Y => n3968);
   U5093 : NOR2X1 port map( A => parameter_A1_div(7), B => n4013, Y => n4011);
   U5094 : NOR2X1 port map( A => parameter_A2_div(7), B => n4056, Y => n4054);
   U5095 : NAND3BX1 port map( AN => n336, B => n339, C => n3695, Y => n3708);
   U5096 : NAND3BX1 port map( AN => n327, B => n330, C => n3743, Y => n3756);
   U5097 : NAND3BX1 port map( AN => n363, B => n366, C => n3791, Y => n3804);
   U5098 : NAND3BX1 port map( AN => n354, B => n357, C => n3839, Y => n3852);
   U5099 : NAND3BX1 port map( AN => n345, B => n348, C => n3647, Y => n3660);
   U5100 : NAND3BX1 port map( AN => parameter_B0_div(7), B => n342, C => n3882,
                           Y => n3895);
   U5101 : NAND3BX1 port map( AN => parameter_B1_div(7), B => n333, C => n3925,
                           Y => n3938);
   U5102 : NAND3BX1 port map( AN => parameter_B2_div(7), B => n324, C => n3968,
                           Y => n3981);
   U5103 : NAND3BX1 port map( AN => parameter_A1_div(7), B => n360, C => n4011,
                           Y => n4024);
   U5104 : NAND3BX1 port map( AN => parameter_A2_div(7), B => n351, C => n4054,
                           Y => n4067);
   U5105 : NOR2BX1 port map( AN => n3705, B => n336, Y => n3704);
   U5106 : NOR2BX1 port map( AN => n3753, B => n327, Y => n3752);
   U5107 : NOR2BX1 port map( AN => n3801, B => n363, Y => n3800);
   U5108 : NOR2BX1 port map( AN => n3849, B => n354, Y => n3848);
   U5109 : NOR2BX1 port map( AN => n3657, B => n345, Y => n3656);
   U5110 : NOR2X1 port map( A => n336, B => n3706, Y => n3705);
   U5111 : NOR2X1 port map( A => n327, B => n3754, Y => n3753);
   U5112 : NOR2X1 port map( A => n363, B => n3802, Y => n3801);
   U5113 : NOR2X1 port map( A => n354, B => n3850, Y => n3849);
   U5114 : NOR2X1 port map( A => n345, B => n3658, Y => n3657);
   U5115 : NOR2BX1 port map( AN => 
                           input_times_b0_div_componentxinput_B_inverted_17_port, B 
                           => n342, Y => 
                           input_times_b0_div_componentxunsigned_B_17);
   U5116 : XOR2X1 port map( A => n3890, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_17_port);
   U5117 : NAND2BX1 port map( AN => parameter_B0_div(7), B => n3891, Y => n3890
                           );
   U5118 : NOR2BX1 port map( AN => 
                           input_p1_times_b1_div_componentxinput_B_inverted_17_port, B 
                           => n333, Y => 
                           input_p1_times_b1_div_componentxunsigned_B_17);
   U5119 : XOR2X1 port map( A => n3933, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_17_port);
   U5120 : NAND2BX1 port map( AN => parameter_B1_div(7), B => n3934, Y => n3933
                           );
   U5121 : NOR2BX1 port map( AN => 
                           input_p2_times_b2_div_componentxinput_B_inverted_17_port, B 
                           => n324, Y => 
                           input_p2_times_b2_div_componentxunsigned_B_17);
   U5122 : XOR2X1 port map( A => n3976, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_17_port);
   U5123 : NAND2BX1 port map( AN => parameter_B2_div(7), B => n3977, Y => n3976
                           );
   U5124 : NOR2BX1 port map( AN => 
                           output_p1_times_a1_div_componentxinput_B_inverted_17_port, B 
                           => n360, Y => 
                           output_p1_times_a1_div_componentxunsigned_B_17);
   U5125 : XOR2X1 port map( A => n4019, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_17_port);
   U5126 : NAND2BX1 port map( AN => parameter_A1_div(7), B => n4020, Y => n4019
                           );
   U5127 : NOR2BX1 port map( AN => 
                           output_p2_times_a2_div_componentxinput_B_inverted_17_port, B 
                           => n351, Y => 
                           output_p2_times_a2_div_componentxunsigned_B_17);
   U5128 : XOR2X1 port map( A => n4062, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_17_port);
   U5129 : NAND2BX1 port map( AN => parameter_A2_div(7), B => n4063, Y => n4062
                           );
   U5130 : OR2X2 port map( A => n3708, B => n336, Y => n3706);
   U5131 : OR2X2 port map( A => n3756, B => n327, Y => n3754);
   U5132 : OR2X2 port map( A => n3804, B => n363, Y => n3802);
   U5133 : OR2X2 port map( A => n3852, B => n354, Y => n3850);
   U5134 : OR2X2 port map( A => n3660, B => n345, Y => n3658);
   U5135 : XOR2X1 port map( A => n847, B => n846, Y => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_1_port);
   U5136 : XOR2X1 port map( A => n1006, B => n1005, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_1_port);
   U5137 : XOR2X1 port map( A => n1165, B => n1164, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_1_port);
   U5138 : XOR2X1 port map( A => n529, B => n528, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_1_port);
   U5139 : XOR2X1 port map( A => n688, B => n687, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_1_port);
   U5140 : XNOR2X1 port map( A => n848, B => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn9, Y 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_2_port);
   U5141 : NOR2X1 port map( A => n846, B => n847, Y => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn9);
   U5142 : XNOR2X1 port map( A => n1007, B => n1765, Y => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_2_port);
   U5143 : NOR2X1 port map( A => n1005, B => n1006, Y => n1765);
   U5144 : XNOR2X1 port map( A => n1166, B => n1774, Y => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_2_port);
   U5145 : NOR2X1 port map( A => n1164, B => n1165, Y => n1774);
   U5146 : XNOR2X1 port map( A => n530, B => n1783, Y => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_2_port);
   U5147 : NOR2X1 port map( A => n528, B => n529, Y => n1783);
   U5148 : XNOR2X1 port map( A => n689, B => n1792, Y => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_2_port);
   U5149 : NOR2X1 port map( A => n687, B => n688, Y => n1792);
   U5150 : INVX1 port map( A => n339, Y => n335);
   U5151 : INVX1 port map( A => n330, Y => n326);
   U5152 : INVX1 port map( A => n366, Y => n362);
   U5153 : INVX1 port map( A => n357, Y => n353);
   U5154 : INVX1 port map( A => n348, Y => n344);
   U5155 : OR3XL port map( A => n847, B => n848, C => n846, Y => 
                           input_times_b0_div_componentxUDxinverter_for_substractionxn8);
   U5156 : OR3XL port map( A => n1006, B => n1007, C => n1005, Y => n1764);
   U5157 : OR3XL port map( A => n1165, B => n1166, C => n1164, Y => n1773);
   U5158 : OR3XL port map( A => n529, B => n530, C => n528, Y => n1782);
   U5159 : OR3XL port map( A => n688, B => n689, C => n687, Y => n1791);
   U5160 : INVX1 port map( A => n342, Y => n341);
   U5161 : INVX1 port map( A => n333, Y => n332);
   U5162 : INVX1 port map( A => n324, Y => n323);
   U5163 : INVX1 port map( A => n360, Y => n359);
   U5164 : INVX1 port map( A => n351, Y => n350);
   U5165 : INVX1 port map( A => n339, Y => n334);
   U5166 : INVX1 port map( A => n330, Y => n325);
   U5167 : INVX1 port map( A => n357, Y => n352);
   U5168 : INVX1 port map( A => n366, Y => n361);
   U5169 : INVX1 port map( A => input_times_b0_div_componentxn48, Y => n849);
   U5170 : INVX1 port map( A => n4226, Y => n1008);
   U5171 : INVX1 port map( A => n4282, Y => n1167);
   U5172 : INVX1 port map( A => n4336, Y => n531);
   U5173 : INVX1 port map( A => n4392, Y => n690);
   U5174 : INVX1 port map( A => input_times_b0_div_componentxn50, Y => n851);
   U5175 : INVX1 port map( A => n4228, Y => n1010);
   U5176 : INVX1 port map( A => n4284, Y => n1169);
   U5177 : INVX1 port map( A => n4338, Y => n533);
   U5178 : INVX1 port map( A => n4394, Y => n692);
   U5179 : INVX1 port map( A => input_times_b0_div_componentxn49, Y => n850);
   U5180 : INVX1 port map( A => n4227, Y => n1009);
   U5181 : INVX1 port map( A => n4283, Y => n1168);
   U5182 : INVX1 port map( A => n4337, Y => n532);
   U5183 : INVX1 port map( A => n4393, Y => n691);
   U5184 : INVX1 port map( A => input_times_b0_div_componentxn51, Y => n852);
   U5185 : INVX1 port map( A => n4229, Y => n1011);
   U5186 : INVX1 port map( A => n4285, Y => n1170);
   U5187 : INVX1 port map( A => n4339, Y => n534);
   U5188 : INVX1 port map( A => n4395, Y => n693);
   U5189 : INVX1 port map( A => input_times_b0_div_componentxn61, Y => n843);
   U5190 : AOI22X1 port map( A0 => n340, A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_16_port, 
                           B1 => n341, Y => input_times_b0_div_componentxn61);
   U5191 : XNOR2X1 port map( A => n3891, B => n340, Y => 
                           input_times_b0_div_componentxinput_B_inverted_16_port);
   U5192 : INVX1 port map( A => n4239, Y => n1002);
   U5193 : AOI22X1 port map( A0 => n331, A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_16_port, 
                           B1 => n332, Y => n4239);
   U5194 : XNOR2X1 port map( A => n3934, B => n331, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_16_port);
   U5195 : INVX1 port map( A => n4295, Y => n1161);
   U5196 : AOI22X1 port map( A0 => n322, A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_16_port, 
                           B1 => n323, Y => n4295);
   U5197 : XNOR2X1 port map( A => n3977, B => n322, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_16_port);
   U5198 : INVX1 port map( A => n4349, Y => n525);
   U5199 : AOI22X1 port map( A0 => n358, A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_16_port, 
                           B1 => n359, Y => n4349);
   U5200 : XNOR2X1 port map( A => n4020, B => n358, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_16_port);
   U5201 : INVX1 port map( A => n4405, Y => n684);
   U5202 : AOI22X1 port map( A0 => n349, A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_16_port, 
                           B1 => n350, Y => n4405);
   U5203 : XNOR2X1 port map( A => n4063, B => n349, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_16_port);
   U5204 : XOR2X1 port map( A => n3703, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_17_port);
   U5205 : NAND2BX1 port map( AN => n336, B => n3704, Y => n3703);
   U5206 : XOR2X1 port map( A => n3751, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_17_port);
   U5207 : NAND2BX1 port map( AN => n327, B => n3752, Y => n3751);
   U5208 : XOR2X1 port map( A => n3847, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_17_port);
   U5209 : NAND2BX1 port map( AN => n354, B => n3848, Y => n3847);
   U5210 : XOR2X1 port map( A => n3655, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_17_port);
   U5211 : NAND2BX1 port map( AN => n345, B => n3656, Y => n3655);
   U5212 : INVX1 port map( A => input_times_b0_div_componentxn47, Y => n848);
   U5213 : INVX1 port map( A => n4225, Y => n1007);
   U5214 : INVX1 port map( A => n4281, Y => n1166);
   U5215 : INVX1 port map( A => n4335, Y => n530);
   U5216 : INVX1 port map( A => n4391, Y => n689);
   U5217 : BUFX3 port map( A => n4409, Y => n172);
   U5218 : AOI22X1 port map( A0 => n335, A1 => n337, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_7_port, 
                           B1 => n335, Y => n4409);
   U5219 : XOR2X1 port map( A => n3697, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_7_port);
   U5220 : BUFX3 port map( A => n4462, Y => n193);
   U5221 : AOI22X1 port map( A0 => n326, A1 => n328, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_7_port, 
                           B1 => n326, Y => n4462);
   U5222 : XOR2X1 port map( A => n3745, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_7_port);
   U5223 : BUFX3 port map( A => n4515, Y => n214);
   U5224 : AOI22X1 port map( A0 => n362, A1 => n364, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_7_port, 
                           B1 => n362, Y => n4515);
   U5225 : XOR2X1 port map( A => n3793, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_7_port);
   U5226 : BUFX3 port map( A => n4568, Y => n235);
   U5227 : AOI22X1 port map( A0 => n353, A1 => n355, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_7_port, 
                           B1 => n353, Y => n4568);
   U5228 : XOR2X1 port map( A => n3841, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_7_port);
   U5229 : BUFX3 port map( A => input_times_b0_mul_componentxn58, Y => n263);
   U5230 : AOI22X1 port map( A0 => n344, A1 => n346, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_7_port
                           , B1 => n344, Y => input_times_b0_mul_componentxn58)
                           ;
   U5231 : XOR2X1 port map( A => n3649, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_7_port
                           );
   U5232 : BUFX3 port map( A => n4408, Y => n171);
   U5233 : AOI22X1 port map( A0 => n334, A1 => n337, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_8_port, 
                           B1 => n335, Y => n4408);
   U5234 : XOR2X1 port map( A => n3696, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_8_port);
   U5235 : OR2X2 port map( A => n336, B => n3697, Y => n3696);
   U5236 : BUFX3 port map( A => n4461, Y => n192);
   U5237 : AOI22X1 port map( A0 => n325, A1 => n328, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_8_port, 
                           B1 => n326, Y => n4461);
   U5238 : XOR2X1 port map( A => n3744, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_8_port);
   U5239 : OR2X2 port map( A => n327, B => n3745, Y => n3744);
   U5240 : BUFX3 port map( A => n4567, Y => n234);
   U5241 : AOI22X1 port map( A0 => n352, A1 => n355, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_8_port, 
                           B1 => n353, Y => n4567);
   U5242 : XOR2X1 port map( A => n3840, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_8_port);
   U5243 : OR2X2 port map( A => n354, B => n3841, Y => n3840);
   U5244 : BUFX3 port map( A => input_times_b0_mul_componentxn57, Y => n262);
   U5245 : AOI22X1 port map( A0 => n344, A1 => n346, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_8_port
                           , B1 => n344, Y => input_times_b0_mul_componentxn57)
                           ;
   U5246 : XOR2X1 port map( A => n3648, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_8_port
                           );
   U5247 : OR2X2 port map( A => n345, B => n3649, Y => n3648);
   U5248 : BUFX3 port map( A => n4514, Y => n213);
   U5249 : AOI22X1 port map( A0 => n361, A1 => n365, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_8_port, 
                           B1 => n362, Y => n4514);
   U5250 : XOR2X1 port map( A => n3792, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_8_port);
   U5251 : OR2X2 port map( A => n363, B => n3793, Y => n3792);
   U5252 : BUFX3 port map( A => n4407, Y => n170);
   U5253 : AOI22X1 port map( A0 => n334, A1 => n337, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_9_port, 
                           B1 => n335, Y => n4407);
   U5254 : XNOR2X1 port map( A => n3695, B => n334, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_9_port);
   U5255 : BUFX3 port map( A => n4460, Y => n191);
   U5256 : AOI22X1 port map( A0 => n325, A1 => n328, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_9_port, 
                           B1 => n326, Y => n4460);
   U5257 : XNOR2X1 port map( A => n3743, B => n325, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_9_port);
   U5258 : BUFX3 port map( A => n4566, Y => n233);
   U5259 : AOI22X1 port map( A0 => n352, A1 => n355, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_9_port, 
                           B1 => n353, Y => n4566);
   U5260 : XNOR2X1 port map( A => n3839, B => n352, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_9_port);
   U5261 : BUFX3 port map( A => input_times_b0_mul_componentxn56, Y => n261);
   U5262 : AOI22X1 port map( A0 => n344, A1 => n346, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_9_port
                           , B1 => n344, Y => input_times_b0_mul_componentxn56)
                           ;
   U5263 : XNOR2X1 port map( A => n3647, B => n343, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_9_port
                           );
   U5264 : BUFX3 port map( A => n4513, Y => n212);
   U5265 : AOI22X1 port map( A0 => n361, A1 => n366, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_9_port, 
                           B1 => n362, Y => n4513);
   U5266 : XNOR2X1 port map( A => n3791, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_9_port);
   U5267 : XOR2X1 port map( A => n3799, B => n361, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_17_port);
   U5268 : NAND2BX1 port map( AN => n363, B => n3800, Y => n3799);
   U5269 : INVX1 port map( A => n283, Y => n317);
   U5270 : INVX1 port map( A => n301, Y => n316);
   U5271 : INVX1 port map( A => n307, Y => n318);
   U5272 : INVX1 port map( A => n308, Y => n315);
   U5273 : BUFX3 port map( A => 
                           output_p2_times_a2_div_componentxoutput_sign_gated, 
                           Y => n169);
   U5274 : BUFX3 port map( A => 
                           output_p1_times_a1_div_componentxoutput_sign_gated, 
                           Y => n168);
   U5275 : BUFX3 port map( A => 
                           input_p1_times_b1_div_componentxoutput_sign_gated, Y
                           => n166);
   U5276 : BUFX3 port map( A => input_times_b0_div_componentxoutput_sign_gated,
                           Y => n260);
   U5277 : INVX1 port map( A => n4359, Y => n1311);
   U5278 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_1, 
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_1_port, 
                           B1 => n169, Y => n4359);
   U5279 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_1, 
                           B => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_0_port, Y 
                           => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_1_port);
   U5280 : INVX1 port map( A => n4193, Y => n1370);
   U5281 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_1, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_1_port, 
                           B1 => n166, Y => n4193);
   U5282 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_1, B
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_0_port, Y 
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_1_port);
   U5283 : OAI2BB1X1 port map( A0N => 
                           output_p1_times_a1_div_componentxUDxshifted_substraction_result_0, 
                           A1N => n371, B0 => n2088, Y => n2108);
   U5284 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_16, 
                           A1 => n2089, B0 => 
                           output_p1_times_a1_div_componentxunsigned_A_17, B1 
                           => n2090, Y => n2088);
   U5285 : NOR2BX1 port map( AN => 
                           output_p1_times_a1_div_componentxinput_A_inverted_17_port, B 
                           => n232, Y => 
                           output_p1_times_a1_div_componentxunsigned_A_17);
   U5286 : XOR2X1 port map( A => n4005, B => n111, Y => 
                           output_p1_times_a1_div_componentxinput_A_inverted_17_port);
   U5287 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_1, 
                           B0 => n2106, Y => n2124);
   U5288 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_0, 
                           A1 => n2089, B0 => n382, B1 => n2090, Y => n2106);
   U5289 : INVX1 port map( A => n4317, Y => n382);
   U5290 : AOI22X1 port map( A0 => n517, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_1_port, 
                           B1 => n112, Y => n4317);
   U5291 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_2, 
                           B0 => n2105, Y => n2123);
   U5292 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_1, 
                           A1 => n2089, B0 => n383, B1 => n2090, Y => n2105);
   U5293 : INVX1 port map( A => n4318, Y => n383);
   U5294 : AOI22X1 port map( A0 => n516, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_2_port, 
                           B1 => n112, Y => n4318);
   U5295 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_3, 
                           B0 => n2104, Y => n2122);
   U5296 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_2, 
                           A1 => n2089, B0 => n384, B1 => n2090, Y => n2104);
   U5297 : INVX1 port map( A => n4319, Y => n384);
   U5298 : AOI22X1 port map( A0 => n509, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_3_port, 
                           B1 => n112, Y => n4319);
   U5299 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_4, 
                           B0 => n2103, Y => n2121);
   U5300 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_3, 
                           A1 => n2089, B0 => n385, B1 => n2090, Y => n2103);
   U5301 : INVX1 port map( A => n4320, Y => n385);
   U5302 : AOI22X1 port map( A0 => n503, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_4_port, 
                           B1 => n112, Y => n4320);
   U5303 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_5, 
                           B0 => n2102, Y => n2120);
   U5304 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_4, 
                           A1 => n2089, B0 => n386, B1 => n2090, Y => n2102);
   U5305 : INVX1 port map( A => n4321, Y => n386);
   U5306 : AOI22X1 port map( A0 => n495, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_5_port, 
                           B1 => n112, Y => n4321);
   U5307 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_6, 
                           B0 => n2101, Y => n2119);
   U5308 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_5, 
                           A1 => n2089, B0 => n387, B1 => n2090, Y => n2101);
   U5309 : INVX1 port map( A => n4322, Y => n387);
   U5310 : AOI22X1 port map( A0 => n488, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_6_port, 
                           B1 => n112, Y => n4322);
   U5311 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_7, 
                           B0 => n2100, Y => n2118);
   U5312 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_6, 
                           A1 => n2089, B0 => n388, B1 => n2090, Y => n2100);
   U5313 : INVX1 port map( A => n4323, Y => n388);
   U5314 : AOI22X1 port map( A0 => n480, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_7_port, 
                           B1 => n112, Y => n4323);
   U5315 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_8, 
                           B0 => n2099, Y => n2117);
   U5316 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_7, 
                           A1 => n2089, B0 => n389, B1 => n2090, Y => n2099);
   U5317 : INVX1 port map( A => n4324, Y => n389);
   U5318 : AOI22X1 port map( A0 => n473, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_8_port, 
                           B1 => n112, Y => n4324);
   U5319 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_9, 
                           B0 => n2098, Y => n2116);
   U5320 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_8, 
                           A1 => n2089, B0 => n390, B1 => n2090, Y => n2098);
   U5321 : INVX1 port map( A => n4325, Y => n390);
   U5322 : AOI22X1 port map( A0 => n463, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_9_port, 
                           B1 => n111, Y => n4325);
   U5323 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_10, 
                           B0 => n2097, Y => n2115);
   U5324 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_9, 
                           A1 => n2089, B0 => n391, B1 => n2090, Y => n2097);
   U5325 : INVX1 port map( A => n4326, Y => n391);
   U5326 : AOI22X1 port map( A0 => n453, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_10_port, 
                           B1 => n111, Y => n4326);
   U5327 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_11, 
                           B0 => n2096, Y => n2114);
   U5328 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_10, 
                           A1 => n2089, B0 => n392, B1 => n2090, Y => n2096);
   U5329 : INVX1 port map( A => n4327, Y => n392);
   U5330 : AOI22X1 port map( A0 => n441, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_11_port, 
                           B1 => n111, Y => n4327);
   U5331 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_12, 
                           B0 => n2095, Y => n2113);
   U5332 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_11, 
                           A1 => n2089, B0 => n393, B1 => n2090, Y => n2095);
   U5333 : INVX1 port map( A => n4328, Y => n393);
   U5334 : AOI22X1 port map( A0 => n432, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_12_port, 
                           B1 => n111, Y => n4328);
   U5335 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_13, 
                           B0 => n2094, Y => n2112);
   U5336 : AOI22XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_12, 
                           A1 => n2089, B0 => n394, B1 => n2090, Y => n2094);
   U5337 : INVX1 port map( A => n4329, Y => n394);
   U5338 : AOI22X1 port map( A0 => n423, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_13_port, 
                           B1 => n111, Y => n4329);
   U5339 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_14, 
                           B0 => n2093, Y => n2111);
   U5340 : AOI22XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_13, 
                           A1 => n2089, B0 => n395, B1 => n2090, Y => n2093);
   U5341 : INVX1 port map( A => n4330, Y => n395);
   U5342 : AOI22X1 port map( A0 => n417, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_14_port, 
                           B1 => n111, Y => n4330);
   U5343 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_15, 
                           B0 => n2092, Y => n2110);
   U5344 : AOI22XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_14, 
                           A1 => n2089, B0 => n396, B1 => n2090, Y => n2092);
   U5345 : INVX1 port map( A => n4331, Y => n396);
   U5346 : AOI22X1 port map( A0 => n408, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_15_port, 
                           B1 => n111, Y => n4331);
   U5347 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_16, 
                           B0 => n2091, Y => n2109);
   U5348 : AOI22XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_15, 
                           A1 => n2089, B0 => n397, B1 => n2090, Y => n2091);
   U5349 : INVX1 port map( A => n4332, Y => n397);
   U5350 : AOI22X1 port map( A0 => n401, A1 => n232, B0 => 
                           output_p1_times_a1_div_componentxinput_A_inverted_16_port, 
                           B1 => n111, Y => n4332);
   U5351 : INVX1 port map( A => n4305, Y => n1331);
   U5352 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_1, 
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_1_port, 
                           B1 => n168, Y => n4305);
   U5353 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_1, 
                           B => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_0_port, Y 
                           => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_1_port);
   U5354 : INVX1 port map( A => input_times_b0_div_componentxn12, Y => n1227);
   U5355 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_1, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_1_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn12);
   U5356 : XOR2X1 port map( A => input_times_b0_div_componentxunsigned_output_1
                           , B => 
                           input_times_b0_div_componentxunsigned_output_inverted_0_port, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_1_port);
   U5357 : NOR3X1 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_7, B
                           => input_p1_times_b1_div_componentxunsigned_output_8
                           , C => n3943, Y => n3941);
   U5358 : NOR3X1 port map( A => input_times_b0_div_componentxunsigned_output_7
                           , B => 
                           input_times_b0_div_componentxunsigned_output_8, C =>
                           n3900, Y => n3898);
   U5359 : NOR3X1 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_7, 
                           B => 
                           output_p2_times_a2_div_componentxunsigned_output_8, 
                           C => n4072, Y => n4070);
   U5360 : NOR3X1 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_7, 
                           B => 
                           output_p1_times_a1_div_componentxunsigned_output_8, 
                           C => n4029, Y => n4027);
   U5361 : INVX1 port map( A => n4303, Y => n1329);
   U5362 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_3, 
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_3_port, 
                           B1 => n168, Y => n4303);
   U5363 : XOR2X1 port map( A => n4033, B => 
                           output_p1_times_a1_div_componentxunsigned_output_3, 
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_3_port);
   U5364 : INVX1 port map( A => input_times_b0_div_componentxn10, Y => n1223);
   U5365 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_3, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_3_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn10);
   U5366 : XOR2X1 port map( A => n3904, B => 
                           input_times_b0_div_componentxunsigned_output_3, Y =>
                           input_times_b0_div_componentxunsigned_output_inverted_3_port);
   U5367 : INVX1 port map( A => n4301, Y => n1327);
   U5368 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_5, 
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_5_port, 
                           B1 => n168, Y => n4301);
   U5369 : XOR2X1 port map( A => n4031, B => 
                           output_p1_times_a1_div_componentxunsigned_output_5, 
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_5_port);
   U5370 : INVX1 port map( A => input_times_b0_div_componentxn8, Y => n1219);
   U5371 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_5, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_5_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn8);
   U5372 : XOR2X1 port map( A => n3902, B => 
                           input_times_b0_div_componentxunsigned_output_5, Y =>
                           input_times_b0_div_componentxunsigned_output_inverted_5_port);
   U5373 : INVX1 port map( A => n4299, Y => n1325);
   U5374 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_7, 
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_7_port, 
                           B1 => n168, Y => n4299);
   U5375 : XOR2X1 port map( A => n4029, B => 
                           output_p1_times_a1_div_componentxunsigned_output_7, 
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_7_port);
   U5376 : INVX1 port map( A => input_times_b0_div_componentxn6, Y => n1215);
   U5377 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_7, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_7_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn6);
   U5378 : XOR2X1 port map( A => n3900, B => 
                           input_times_b0_div_componentxunsigned_output_7, Y =>
                           input_times_b0_div_componentxunsigned_output_inverted_7_port);
   U5379 : INVX1 port map( A => n4201, Y => n1378);
   U5380 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_10, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_10_port, 
                           B1 => n166, Y => n4201);
   U5381 : XOR2X1 port map( A => n3956, B => 
                           input_p1_times_b1_div_componentxunsigned_output_10, 
                           Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_10_port);
   U5382 : NAND2X1 port map( A => n3941, B => n1448, Y => n3956);
   U5383 : INVX1 port map( A => input_times_b0_div_componentxn17, Y => n1232);
   U5384 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_13, A1 
                           => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_13_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn17);
   U5385 : XOR2X1 port map( A => n3909, B => 
                           input_times_b0_div_componentxunsigned_output_13, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_13_port);
   U5386 : NAND3BX1 port map( AN => 
                           input_p1_times_b1_div_componentxunsigned_output_10, 
                           B => n1448, C => n3941, Y => n3954);
   U5387 : NAND3BX1 port map( AN => 
                           input_times_b0_div_componentxunsigned_output_10, B 
                           => n1272, C => n3898, Y => n3911);
   U5388 : OR3XL port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_5, 
                           B => 
                           output_p2_times_a2_div_componentxunsigned_output_6, 
                           C => n4074, Y => n4072);
   U5389 : OR3XL port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_5, 
                           B => 
                           output_p1_times_a1_div_componentxunsigned_output_6, 
                           C => n4031, Y => n4029);
   U5390 : OR3XL port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_5, B
                           => input_p1_times_b1_div_componentxunsigned_output_6
                           , C => n3945, Y => n3943);
   U5391 : OR3XL port map( A => input_times_b0_div_componentxunsigned_output_5,
                           B => input_times_b0_div_componentxunsigned_output_6,
                           C => n3902, Y => n3900);
   U5392 : OR3XL port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_11, 
                           B => 
                           input_p1_times_b1_div_componentxunsigned_output_12, 
                           C => n3954, Y => n3952);
   U5393 : OR3XL port map( A => input_times_b0_div_componentxunsigned_output_11
                           , B => 
                           input_times_b0_div_componentxunsigned_output_12, C 
                           => n3911, Y => n3909);
   U5394 : BUFX3 port map( A => 
                           input_p2_times_b2_div_componentxoutput_sign_gated, Y
                           => n167);
   U5395 : OR3XL port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_1, 
                           B => 
                           output_p2_times_a2_div_componentxunsigned_output_2, 
                           C => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_0_port, Y 
                           => n4076);
   U5396 : OR3XL port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_1, 
                           B => 
                           output_p1_times_a1_div_componentxunsigned_output_2, 
                           C => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_0_port, Y 
                           => n4033);
   U5397 : OR3XL port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_1, B
                           => input_p1_times_b1_div_componentxunsigned_output_2
                           , C => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_0_port, Y 
                           => n3947);
   U5398 : OR3XL port map( A => input_times_b0_div_componentxunsigned_output_1,
                           B => input_times_b0_div_componentxunsigned_output_2,
                           C => 
                           input_times_b0_div_componentxunsigned_output_inverted_0_port, Y 
                           => n3904);
   U5399 : OR3XL port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_1, B
                           => input_p2_times_b2_div_componentxunsigned_output_2
                           , C => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_0_port, Y 
                           => n3990);
   U5400 : OR3XL port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_3, 
                           B => 
                           output_p2_times_a2_div_componentxunsigned_output_4, 
                           C => n4076, Y => n4074);
   U5401 : OR3XL port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_3, 
                           B => 
                           output_p1_times_a1_div_componentxunsigned_output_4, 
                           C => n4033, Y => n4031);
   U5402 : OR3XL port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_3, B
                           => input_p1_times_b1_div_componentxunsigned_output_4
                           , C => n3947, Y => n3945);
   U5403 : OR3XL port map( A => input_times_b0_div_componentxunsigned_output_3,
                           B => input_times_b0_div_componentxunsigned_output_4,
                           C => n3904, Y => n3902);
   U5404 : INVX1 port map( A => input_times_b0_div_componentxn21, Y => n1237);
   U5405 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_0_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn21);
   U5406 : INVX1 port map( A => n4314, Y => n1340);
   U5407 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_0_port, 
                           B1 => n168, Y => n4314);
   U5408 : INVX1 port map( A => n4357, Y => n1309);
   U5409 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_3, 
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_3_port, 
                           B1 => n169, Y => n4357);
   U5410 : XOR2X1 port map( A => n4076, B => 
                           output_p2_times_a2_div_componentxunsigned_output_3, 
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_3_port);
   U5411 : INVX1 port map( A => n4191, Y => n1368);
   U5412 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_3, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_3_port, 
                           B1 => n166, Y => n4191);
   U5413 : XOR2X1 port map( A => n3947, B => 
                           input_p1_times_b1_div_componentxunsigned_output_3, Y
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_3_port);
   U5414 : INVX1 port map( A => n4355, Y => n1307);
   U5415 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_5, 
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_5_port, 
                           B1 => n169, Y => n4355);
   U5416 : XOR2X1 port map( A => n4074, B => 
                           output_p2_times_a2_div_componentxunsigned_output_5, 
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_5_port);
   U5417 : INVX1 port map( A => n4247, Y => n1348);
   U5418 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_3, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_3_port, 
                           B1 => n167, Y => n4247);
   U5419 : XOR2X1 port map( A => n3990, B => 
                           input_p2_times_b2_div_componentxunsigned_output_3, Y
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_3_port);
   U5420 : INVX1 port map( A => n4189, Y => n1366);
   U5421 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_5, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_5_port, 
                           B1 => n166, Y => n4189);
   U5422 : XOR2X1 port map( A => n3945, B => 
                           input_p1_times_b1_div_componentxunsigned_output_5, Y
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_5_port);
   U5423 : INVX1 port map( A => n4353, Y => n1305);
   U5424 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_7, 
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_7_port, 
                           B1 => n169, Y => n4353);
   U5425 : XOR2X1 port map( A => n4072, B => 
                           output_p2_times_a2_div_componentxunsigned_output_7, 
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_7_port);
   U5426 : INVX1 port map( A => n4187, Y => n1364);
   U5427 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_7, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_7_port, 
                           B1 => n166, Y => n4187);
   U5428 : XOR2X1 port map( A => n3943, B => 
                           input_p1_times_b1_div_componentxunsigned_output_7, Y
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_7_port);
   U5429 : INVX1 port map( A => n4351, Y => n1303);
   U5430 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_9, 
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_9_port, 
                           B1 => n169, Y => n4351);
   U5431 : XNOR2X1 port map( A => n4070, B => 
                           output_p2_times_a2_div_componentxunsigned_output_9, 
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_9_port);
   U5432 : INVX1 port map( A => n4185, Y => n1362);
   U5433 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_9, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_9_port, 
                           B1 => n166, Y => n4185);
   U5434 : XNOR2X1 port map( A => n3941, B => 
                           input_p1_times_b1_div_componentxunsigned_output_9, Y
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_9_port);
   U5435 : INVX1 port map( A => n4198, Y => n1375);
   U5436 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_13, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_13_port, 
                           B1 => n166, Y => n4198);
   U5437 : XOR2X1 port map( A => n3952, B => 
                           input_p1_times_b1_div_componentxunsigned_output_13, 
                           Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_13_port);
   U5438 : INVX1 port map( A => n4202, Y => n1379);
   U5439 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_0_port, 
                           B1 => n166, Y => n4202);
   U5440 : INVX1 port map( A => n4368, Y => n1320);
   U5441 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_0_port, 
                           B1 => n169, Y => n4368);
   U5442 : INVX1 port map( A => n4258, Y => n1359);
   U5443 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_0_port, 
                           B1 => n167, Y => n4258);
   U5444 : INVX1 port map( A => n4200, Y => n1377);
   U5445 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_11, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_11_port, 
                           B1 => n166, Y => n4200);
   U5446 : XOR2X1 port map( A => n3954, B => 
                           input_p1_times_b1_div_componentxunsigned_output_11, 
                           Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_11_port);
   U5447 : INVX1 port map( A => input_times_b0_div_componentxn19, Y => n1234);
   U5448 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_11, A1 
                           => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_11_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn19);
   U5449 : XOR2X1 port map( A => n3911, B => 
                           input_times_b0_div_componentxunsigned_output_11, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_11_port);
   U5450 : INVX1 port map( A => n4249, Y => n1350);
   U5451 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_1, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_1_port, 
                           B1 => n167, Y => n4249);
   U5452 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_1, B
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_0_port, Y 
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_1_port);
   U5453 : INVX1 port map( A => n4297, Y => n1323);
   U5454 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_9, 
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_9_port, 
                           B1 => n168, Y => n4297);
   U5455 : XNOR2X1 port map( A => n4027, B => 
                           output_p1_times_a1_div_componentxunsigned_output_9, 
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_9_port);
   U5456 : INVX1 port map( A => input_times_b0_div_componentxn3, Y => n1211);
   U5457 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_9, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_9_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn3);
   U5458 : XNOR2X1 port map( A => n3898, B => 
                           input_times_b0_div_componentxunsigned_output_9, Y =>
                           input_times_b0_div_componentxunsigned_output_inverted_9_port);
   U5459 : INVX1 port map( A => n4358, Y => n1310);
   U5460 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_2, 
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_2_port, 
                           B1 => n169, Y => n4358);
   U5461 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_2, 
                           B => n4077, Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_2_port);
   U5462 : NOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_0_port, B 
                           => 
                           output_p2_times_a2_div_componentxunsigned_output_1, 
                           Y => n4077);
   U5463 : INVX1 port map( A => n4192, Y => n1369);
   U5464 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_2, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_2_port, 
                           B1 => n166, Y => n4192);
   U5465 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_2, B
                           => n3948, Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_2_port);
   U5466 : NOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_0_port, B 
                           => input_p1_times_b1_div_componentxunsigned_output_1
                           , Y => n3948);
   U5467 : INVX1 port map( A => n4356, Y => n1308);
   U5468 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_4, 
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_4_port, 
                           B1 => n169, Y => n4356);
   U5469 : XOR2X1 port map( A => n4075, B => 
                           output_p2_times_a2_div_componentxunsigned_output_4, 
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_4_port);
   U5470 : OR2X2 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_3, 
                           B => n4076, Y => n4075);
   U5471 : INVX1 port map( A => n4248, Y => n1349);
   U5472 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_2, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_2_port, 
                           B1 => n167, Y => n4248);
   U5473 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_2, B
                           => n3991, Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_2_port);
   U5474 : NOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_0_port, B 
                           => input_p2_times_b2_div_componentxunsigned_output_1
                           , Y => n3991);
   U5475 : INVX1 port map( A => n4190, Y => n1367);
   U5476 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_4, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_4_port, 
                           B1 => n166, Y => n4190);
   U5477 : XOR2X1 port map( A => n3946, B => 
                           input_p1_times_b1_div_componentxunsigned_output_4, Y
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_4_port);
   U5478 : OR2X2 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_3, B
                           => n3947, Y => n3946);
   U5479 : INVX1 port map( A => n4354, Y => n1306);
   U5480 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_6, 
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_6_port, 
                           B1 => n169, Y => n4354);
   U5481 : XOR2X1 port map( A => n4073, B => 
                           output_p2_times_a2_div_componentxunsigned_output_6, 
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_6_port);
   U5482 : OR2X2 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_5, 
                           B => n4074, Y => n4073);
   U5483 : INVX1 port map( A => n4188, Y => n1365);
   U5484 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_6, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_6_port, 
                           B1 => n166, Y => n4188);
   U5485 : XOR2X1 port map( A => n3944, B => 
                           input_p1_times_b1_div_componentxunsigned_output_6, Y
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_6_port);
   U5486 : OR2X2 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_5, B
                           => n3945, Y => n3944);
   U5487 : INVX1 port map( A => n4352, Y => n1304);
   U5488 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_8, 
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_8_port, 
                           B1 => n169, Y => n4352);
   U5489 : XOR2X1 port map( A => n4071, B => 
                           output_p2_times_a2_div_componentxunsigned_output_8, 
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_8_port);
   U5490 : OR2X2 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_7, 
                           B => n4072, Y => n4071);
   U5491 : INVX1 port map( A => n4186, Y => n1363);
   U5492 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_8, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_8_port, 
                           B1 => n166, Y => n4186);
   U5493 : XOR2X1 port map( A => n3942, B => 
                           input_p1_times_b1_div_componentxunsigned_output_8, Y
                           => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_8_port);
   U5494 : OR2X2 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_7, B
                           => n3943, Y => n3942);
   U5495 : INVX1 port map( A => n4199, Y => n1376);
   U5496 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_12, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_12_port, 
                           B1 => n166, Y => n4199);
   U5497 : XOR2X1 port map( A => n3955, B => 
                           input_p1_times_b1_div_componentxunsigned_output_12, 
                           Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_12_port);
   U5498 : OR2X2 port map( A => n3954, B => 
                           input_p1_times_b1_div_componentxunsigned_output_11, 
                           Y => n3955);
   U5499 : INVX1 port map( A => n4197, Y => n1374);
   U5500 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_14, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_14_port, 
                           B1 => n166, Y => n4197);
   U5501 : XOR2X1 port map( A => n3953, B => 
                           input_p1_times_b1_div_componentxunsigned_output_14, 
                           Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_14_port);
   U5502 : OR2X2 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_13, 
                           B => n3952, Y => n3953);
   U5503 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxinput_containerxparallel_out_0, 
                           B0 => n2107, Y => n2125);
   U5504 : NAND2XL port map( A => n381, B => n2090, Y => n2107);
   U5505 : INVX1 port map( A => n4316, Y => n381);
   U5506 : AOI22X1 port map( A0 => n518, A1 => n232, B0 => n518, B1 => n112, Y 
                           => n4316);
   U5507 : INVX1 port map( A => n4304, Y => n1330);
   U5508 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_2, 
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_2_port, 
                           B1 => n168, Y => n4304);
   U5509 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_2, 
                           B => n4034, Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_2_port);
   U5510 : NOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_0_port, B 
                           => 
                           output_p1_times_a1_div_componentxunsigned_output_1, 
                           Y => n4034);
   U5511 : INVX1 port map( A => input_times_b0_div_componentxn11, Y => n1225);
   U5512 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_2, A1 
                           => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_2_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn11);
   U5513 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxunsigned_output_2, B =>
                           n3905, Y => 
                           input_times_b0_div_componentxunsigned_output_inverted_2_port);
   U5514 : NOR2X1 port map( A => 
                           input_times_b0_div_componentxunsigned_output_inverted_0_port, B 
                           => input_times_b0_div_componentxunsigned_output_1, Y
                           => n3905);
   U5515 : INVX1 port map( A => n4302, Y => n1328);
   U5516 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_4, 
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_4_port, 
                           B1 => n168, Y => n4302);
   U5517 : XOR2X1 port map( A => n4032, B => 
                           output_p1_times_a1_div_componentxunsigned_output_4, 
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_4_port);
   U5518 : OR2X2 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_3, 
                           B => n4033, Y => n4032);
   U5519 : INVX1 port map( A => input_times_b0_div_componentxn9, Y => n1221);
   U5520 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_4, A1 
                           => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_4_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn9);
   U5521 : XOR2X1 port map( A => n3903, B => 
                           input_times_b0_div_componentxunsigned_output_4, Y =>
                           input_times_b0_div_componentxunsigned_output_inverted_4_port);
   U5522 : OR2X2 port map( A => input_times_b0_div_componentxunsigned_output_3,
                           B => n3904, Y => n3903);
   U5523 : INVX1 port map( A => n4300, Y => n1326);
   U5524 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_6, 
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_6_port, 
                           B1 => n168, Y => n4300);
   U5525 : XOR2X1 port map( A => n4030, B => 
                           output_p1_times_a1_div_componentxunsigned_output_6, 
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_6_port);
   U5526 : OR2X2 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_5, 
                           B => n4031, Y => n4030);
   U5527 : INVX1 port map( A => input_times_b0_div_componentxn7, Y => n1217);
   U5528 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_6, A1 
                           => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_6_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn7);
   U5529 : XOR2X1 port map( A => n3901, B => 
                           input_times_b0_div_componentxunsigned_output_6, Y =>
                           input_times_b0_div_componentxunsigned_output_inverted_6_port);
   U5530 : OR2X2 port map( A => input_times_b0_div_componentxunsigned_output_5,
                           B => n3902, Y => n3901);
   U5531 : INVX1 port map( A => n4298, Y => n1324);
   U5532 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_8, 
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_8_port, 
                           B1 => n168, Y => n4298);
   U5533 : XOR2X1 port map( A => n4028, B => 
                           output_p1_times_a1_div_componentxunsigned_output_8, 
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_8_port);
   U5534 : OR2X2 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_7, 
                           B => n4029, Y => n4028);
   U5535 : INVX1 port map( A => input_times_b0_div_componentxn5, Y => n1213);
   U5536 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_8, A1 
                           => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_8_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn5);
   U5537 : XOR2X1 port map( A => n3899, B => 
                           input_times_b0_div_componentxunsigned_output_8, Y =>
                           input_times_b0_div_componentxunsigned_output_inverted_8_port);
   U5538 : OR2X2 port map( A => input_times_b0_div_componentxunsigned_output_7,
                           B => n3900, Y => n3899);
   U5539 : INVX1 port map( A => input_times_b0_div_componentxn20, Y => n1235);
   U5540 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_10, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_10_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn20);
   U5541 : XOR2X1 port map( A => n3913, B => 
                           input_times_b0_div_componentxunsigned_output_10, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_10_port);
   U5542 : NAND2X1 port map( A => n3898, B => n1272, Y => n3913);
   U5543 : INVX1 port map( A => input_times_b0_div_componentxn18, Y => n1233);
   U5544 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_12, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_12_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn18);
   U5545 : XOR2X1 port map( A => n3912, B => 
                           input_times_b0_div_componentxunsigned_output_12, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_12_port);
   U5546 : OR2X2 port map( A => n3911, B => 
                           input_times_b0_div_componentxunsigned_output_11, Y 
                           => n3912);
   U5547 : OAI2BB2X1 port map( B0 => n108, B1 => n147, A0N => n4315, A1N => 
                           n108, Y => n4350);
   U5548 : AND2X2 port map( A => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , B => en, Y => n108);
   U5549 : NOR3X1 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_7, B
                           => input_p2_times_b2_div_componentxunsigned_output_8
                           , C => n3986, Y => n3984);
   U5550 : NOR3X1 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_13, 
                           B => 
                           input_p1_times_b1_div_componentxunsigned_output_14, 
                           C => n3952, Y => n3951);
   U5551 : NOR3X1 port map( A => 
                           input_times_b0_div_componentxunsigned_output_13, B 
                           => input_times_b0_div_componentxunsigned_output_14, 
                           C => n3909, Y => n3908);
   U5552 : NOR3X1 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_13,
                           B => 
                           output_p2_times_a2_div_componentxunsigned_output_14,
                           C => n4081, Y => n4080);
   U5553 : NOR3X1 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_13,
                           B => 
                           output_p1_times_a1_div_componentxunsigned_output_14,
                           C => n4038, Y => n4037);
   U5554 : NOR3X1 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_13, 
                           B => 
                           input_p2_times_b2_div_componentxunsigned_output_14, 
                           C => n3995, Y => n3994);
   U5555 : INVX1 port map( A => n4367, Y => n1319);
   U5556 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_10,
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_10_port, 
                           B1 => n169, Y => n4367);
   U5557 : XOR2X1 port map( A => n4085, B => 
                           output_p2_times_a2_div_componentxunsigned_output_10,
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_10_port);
   U5558 : NAND2X1 port map( A => n4070, B => n1391, Y => n4085);
   U5559 : INVX1 port map( A => n4257, Y => n1358);
   U5560 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_10, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_10_port, 
                           B1 => n167, Y => n4257);
   U5561 : XOR2X1 port map( A => n3999, B => 
                           input_p2_times_b2_div_componentxunsigned_output_10, 
                           Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_10_port);
   U5562 : NAND2X1 port map( A => n3984, B => n1429, Y => n3999);
   U5563 : INVX1 port map( A => n4310, Y => n1336);
   U5564 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_13,
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_13_port, 
                           B1 => n168, Y => n4310);
   U5565 : XOR2X1 port map( A => n4038, B => 
                           output_p1_times_a1_div_componentxunsigned_output_13,
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_13_port);
   U5566 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_17, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_17_port, 
                           B1 => n166, Y => n4194);
   U5567 : XOR2X1 port map( A => n3949, B => 
                           input_p1_times_b1_div_componentxunsigned_output_17, 
                           Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_17_port);
   U5568 : NAND2BX1 port map( AN => 
                           input_p1_times_b1_div_componentxunsigned_output_16, 
                           B => n3950, Y => n3949);
   U5569 : NAND3BX1 port map( AN => 
                           output_p2_times_a2_div_componentxunsigned_output_10,
                           B => n1391, C => n4070, Y => n4083);
   U5570 : NAND3BX1 port map( AN => 
                           output_p1_times_a1_div_componentxunsigned_output_10,
                           B => n1410, C => n4027, Y => n4040);
   U5571 : NAND3BX1 port map( AN => 
                           input_p2_times_b2_div_componentxunsigned_output_10, 
                           B => n1429, C => n3984, Y => n3997);
   U5572 : NOR2BX1 port map( AN => n3951, B => 
                           input_p1_times_b1_div_componentxunsigned_output_15, 
                           Y => n3950);
   U5573 : NOR2BX1 port map( AN => n3908, B => 
                           input_times_b0_div_componentxunsigned_output_15, Y 
                           => n3907);
   U5574 : NOR2BX1 port map( AN => n4037, B => 
                           output_p1_times_a1_div_componentxunsigned_output_15,
                           Y => n4036);
   U5575 : NOR2BX1 port map( AN => n4080, B => 
                           output_p2_times_a2_div_componentxunsigned_output_15,
                           Y => n4079);
   U5576 : NOR2BX1 port map( AN => n3994, B => 
                           input_p2_times_b2_div_componentxunsigned_output_15, 
                           Y => n3993);
   U5577 : OR3XL port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_5, B
                           => input_p2_times_b2_div_componentxunsigned_output_6
                           , C => n3988, Y => n3986);
   U5578 : OR3XL port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_11,
                           B => 
                           output_p2_times_a2_div_componentxunsigned_output_12,
                           C => n4083, Y => n4081);
   U5579 : OR3XL port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_11,
                           B => 
                           output_p1_times_a1_div_componentxunsigned_output_12,
                           C => n4040, Y => n4038);
   U5580 : OR3XL port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_11, 
                           B => 
                           input_p2_times_b2_div_componentxunsigned_output_12, 
                           C => n3997, Y => n3995);
   U5581 : OR3XL port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_3, B
                           => input_p2_times_b2_div_componentxunsigned_output_4
                           , C => n3990, Y => n3988);
   U5582 : INVX1 port map( A => n4245, Y => n1346);
   U5583 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_5, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_5_port, 
                           B1 => n167, Y => n4245);
   U5584 : XOR2X1 port map( A => n3988, B => 
                           input_p2_times_b2_div_componentxunsigned_output_5, Y
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_5_port);
   U5585 : INVX1 port map( A => n4243, Y => n1344);
   U5586 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_7, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_7_port, 
                           B1 => n167, Y => n4243);
   U5587 : XOR2X1 port map( A => n3986, B => 
                           input_p2_times_b2_div_componentxunsigned_output_7, Y
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_7_port);
   U5588 : INVX1 port map( A => n4241, Y => n1342);
   U5589 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_9, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_9_port, 
                           B1 => n167, Y => n4241);
   U5590 : XNOR2X1 port map( A => n3984, B => 
                           input_p2_times_b2_div_componentxunsigned_output_9, Y
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_9_port);
   U5591 : INVX1 port map( A => n4364, Y => n1316);
   U5592 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_13,
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_13_port, 
                           B1 => n169, Y => n4364);
   U5593 : XOR2X1 port map( A => n4081, B => 
                           output_p2_times_a2_div_componentxunsigned_output_13,
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_13_port);
   U5594 : INVX1 port map( A => n4254, Y => n1355);
   U5595 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_13, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_13_port, 
                           B1 => n167, Y => n4254);
   U5596 : XOR2X1 port map( A => n3995, B => 
                           input_p2_times_b2_div_componentxunsigned_output_13, 
                           Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_13_port);
   U5597 : INVX1 port map( A => n4196, Y => n1373);
   U5598 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_15, 
                           A1 => n151, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_15_port, 
                           B1 => n166, Y => n4196);
   U5599 : XNOR2X1 port map( A => n3951, B => 
                           input_p1_times_b1_div_componentxunsigned_output_15, 
                           Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_15_port);
   U5600 : INVX1 port map( A => n4362, Y => n1314);
   U5601 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_15,
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_15_port, 
                           B1 => n169, Y => n4362);
   U5602 : XNOR2X1 port map( A => n4080, B => 
                           output_p2_times_a2_div_componentxunsigned_output_15,
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_15_port);
   U5603 : INVX1 port map( A => n4252, Y => n1353);
   U5604 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_15, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_15_port, 
                           B1 => n167, Y => n4252);
   U5605 : XNOR2X1 port map( A => n3994, B => 
                           input_p2_times_b2_div_componentxunsigned_output_15, 
                           Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_15_port);
   U5606 : INVX1 port map( A => n4195, Y => n1372);
   U5607 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_16, 
                           A1 => n152, B0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_16_port, 
                           B1 => n166, Y => n4195);
   U5608 : XNOR2X1 port map( A => n3950, B => 
                           input_p1_times_b1_div_componentxunsigned_output_16, 
                           Y => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_16_port);
   U5609 : INVX1 port map( A => n4361, Y => n1313);
   U5610 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_16,
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_16_port, 
                           B1 => n169, Y => n4361);
   U5611 : XNOR2X1 port map( A => n4079, B => 
                           output_p2_times_a2_div_componentxunsigned_output_16,
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_16_port);
   U5612 : INVX1 port map( A => n4251, Y => n1352);
   U5613 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_16, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_16_port, 
                           B1 => n167, Y => n4251);
   U5614 : XNOR2X1 port map( A => n3993, B => 
                           input_p2_times_b2_div_componentxunsigned_output_16, 
                           Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_16_port);
   U5615 : INVX1 port map( A => n4366, Y => n1318);
   U5616 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_11,
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_11_port, 
                           B1 => n169, Y => n4366);
   U5617 : XOR2X1 port map( A => n4083, B => 
                           output_p2_times_a2_div_componentxunsigned_output_11,
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_11_port);
   U5618 : INVX1 port map( A => n4312, Y => n1338);
   U5619 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_11,
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_11_port, 
                           B1 => n168, Y => n4312);
   U5620 : XOR2X1 port map( A => n4040, B => 
                           output_p1_times_a1_div_componentxunsigned_output_11,
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_11_port);
   U5621 : INVX1 port map( A => n4256, Y => n1357);
   U5622 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_11, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_11_port, 
                           B1 => n167, Y => n4256);
   U5623 : XOR2X1 port map( A => n3997, B => 
                           input_p2_times_b2_div_componentxunsigned_output_11, 
                           Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_11_port);
   U5624 : INVX1 port map( A => input_times_b0_div_componentxn15, Y => n1230);
   U5625 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_15, A1 
                           => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_15_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn15);
   U5626 : XNOR2X1 port map( A => n3908, B => 
                           input_times_b0_div_componentxunsigned_output_15, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_15_port);
   U5627 : INVX1 port map( A => n4308, Y => n1334);
   U5628 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_15,
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_15_port, 
                           B1 => n168, Y => n4308);
   U5629 : XNOR2X1 port map( A => n4037, B => 
                           output_p1_times_a1_div_componentxunsigned_output_15,
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_15_port);
   U5630 : INVX1 port map( A => n4246, Y => n1347);
   U5631 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_4, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_4_port, 
                           B1 => n167, Y => n4246);
   U5632 : XOR2X1 port map( A => n3989, B => 
                           input_p2_times_b2_div_componentxunsigned_output_4, Y
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_4_port);
   U5633 : OR2X2 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_3, B
                           => n3990, Y => n3989);
   U5634 : INVX1 port map( A => n4244, Y => n1345);
   U5635 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_6, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_6_port, 
                           B1 => n167, Y => n4244);
   U5636 : XOR2X1 port map( A => n3987, B => 
                           input_p2_times_b2_div_componentxunsigned_output_6, Y
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_6_port);
   U5637 : OR2X2 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_5, B
                           => n3988, Y => n3987);
   U5638 : INVX1 port map( A => n4242, Y => n1343);
   U5639 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_8, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_8_port, 
                           B1 => n167, Y => n4242);
   U5640 : XOR2X1 port map( A => n3985, B => 
                           input_p2_times_b2_div_componentxunsigned_output_8, Y
                           => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_8_port);
   U5641 : OR2X2 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_7, B
                           => n3986, Y => n3985);
   U5642 : INVX1 port map( A => n4365, Y => n1317);
   U5643 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_12,
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_12_port, 
                           B1 => n169, Y => n4365);
   U5644 : XOR2X1 port map( A => n4084, B => 
                           output_p2_times_a2_div_componentxunsigned_output_12,
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_12_port);
   U5645 : OR2X2 port map( A => n4083, B => 
                           output_p2_times_a2_div_componentxunsigned_output_11,
                           Y => n4084);
   U5646 : INVX1 port map( A => n4255, Y => n1356);
   U5647 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_12, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_12_port, 
                           B1 => n167, Y => n4255);
   U5648 : XOR2X1 port map( A => n3998, B => 
                           input_p2_times_b2_div_componentxunsigned_output_12, 
                           Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_12_port);
   U5649 : OR2X2 port map( A => n3997, B => 
                           input_p2_times_b2_div_componentxunsigned_output_11, 
                           Y => n3998);
   U5650 : INVX1 port map( A => n4363, Y => n1315);
   U5651 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_14,
                           A1 => n146, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_14_port, 
                           B1 => n169, Y => n4363);
   U5652 : XOR2X1 port map( A => n4082, B => 
                           output_p2_times_a2_div_componentxunsigned_output_14,
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_14_port);
   U5653 : OR2X2 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_13,
                           B => n4081, Y => n4082);
   U5654 : INVX1 port map( A => n4253, Y => n1354);
   U5655 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_14, 
                           A1 => n150, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_14_port, 
                           B1 => n167, Y => n4253);
   U5656 : XOR2X1 port map( A => n3996, B => 
                           input_p2_times_b2_div_componentxunsigned_output_14, 
                           Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_14_port);
   U5657 : OR2X2 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_13, 
                           B => n3995, Y => n3996);
   U5658 : INVX1 port map( A => input_times_b0_div_componentxn14, Y => n1229);
   U5659 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_16, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_16_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn14);
   U5660 : XNOR2X1 port map( A => n3907, B => 
                           input_times_b0_div_componentxunsigned_output_16, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_16_port);
   U5661 : INVX1 port map( A => n4307, Y => n1333);
   U5662 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_16,
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_16_port, 
                           B1 => n168, Y => n4307);
   U5663 : XNOR2X1 port map( A => n4036, B => 
                           output_p1_times_a1_div_componentxunsigned_output_16,
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_16_port);
   U5664 : INVX1 port map( A => n4313, Y => n1339);
   U5665 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_10,
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_10_port, 
                           B1 => n168, Y => n4313);
   U5666 : XOR2X1 port map( A => n4042, B => 
                           output_p1_times_a1_div_componentxunsigned_output_10,
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_10_port);
   U5667 : NAND2X1 port map( A => n4027, B => n1410, Y => n4042);
   U5668 : INVX1 port map( A => n4311, Y => n1337);
   U5669 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_12,
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_12_port, 
                           B1 => n168, Y => n4311);
   U5670 : XOR2X1 port map( A => n4041, B => 
                           output_p1_times_a1_div_componentxunsigned_output_12,
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_12_port);
   U5671 : OR2X2 port map( A => n4040, B => 
                           output_p1_times_a1_div_componentxunsigned_output_11,
                           Y => n4041);
   U5672 : INVX1 port map( A => input_times_b0_div_componentxn16, Y => n1231);
   U5673 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_14, A1 
                           => n136, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_14_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn16);
   U5674 : XOR2X1 port map( A => n3910, B => 
                           input_times_b0_div_componentxunsigned_output_14, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_14_port);
   U5675 : OR2X2 port map( A => input_times_b0_div_componentxunsigned_output_13
                           , B => n3909, Y => n3910);
   U5676 : INVX1 port map( A => n4309, Y => n1335);
   U5677 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_14,
                           A1 => n148, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_14_port, 
                           B1 => n168, Y => n4309);
   U5678 : XOR2X1 port map( A => n4039, B => 
                           output_p1_times_a1_div_componentxunsigned_output_14,
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_14_port);
   U5679 : OR2X2 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_13,
                           B => n4038, Y => n4039);
   U5680 : INVX1 port map( A => input_times_b0_div_componentxn13, Y => n1228);
   U5681 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_17, A1 
                           => n135, B0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_17_port, 
                           B1 => n260, Y => input_times_b0_div_componentxn13);
   U5682 : XOR2X1 port map( A => n3906, B => 
                           input_times_b0_div_componentxunsigned_output_17, Y 
                           => 
                           input_times_b0_div_componentxunsigned_output_inverted_17_port);
   U5683 : NAND2BX1 port map( AN => 
                           input_times_b0_div_componentxunsigned_output_16, B 
                           => n3907, Y => n3906);
   U5684 : INVX1 port map( A => n4306, Y => n1332);
   U5685 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_17,
                           A1 => n147, B0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_17_port, 
                           B1 => n168, Y => n4306);
   U5686 : XOR2X1 port map( A => n4035, B => 
                           output_p1_times_a1_div_componentxunsigned_output_17,
                           Y => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_17_port);
   U5687 : NAND2BX1 port map( AN => 
                           output_p1_times_a1_div_componentxunsigned_output_16,
                           B => n4036, Y => n4035);
   U5688 : INVX1 port map( A => n4360, Y => n1312);
   U5689 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_17,
                           A1 => n145, B0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_17_port, 
                           B1 => n169, Y => n4360);
   U5690 : XOR2X1 port map( A => n4078, B => 
                           output_p2_times_a2_div_componentxunsigned_output_17,
                           Y => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_17_port);
   U5691 : NAND2BX1 port map( AN => 
                           output_p2_times_a2_div_componentxunsigned_output_16,
                           B => n4079, Y => n4078);
   U5692 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_17, 
                           A1 => n149, B0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_17_port, 
                           B1 => n167, Y => n4250);
   U5693 : XOR2X1 port map( A => n3992, B => 
                           input_p2_times_b2_div_componentxunsigned_output_17, 
                           Y => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_17_port);
   U5694 : NAND2BX1 port map( AN => 
                           input_p2_times_b2_div_componentxunsigned_output_16, 
                           B => n3993, Y => n3992);
   U5695 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxunsigned_output_9, Y
                           => n1448);
   U5696 : INVX1 port map( A => input_times_b0_div_componentxunsigned_output_9,
                           Y => n1272);
   U5697 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxunsigned_output_9, 
                           Y => n1391);
   U5698 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxunsigned_output_9, 
                           Y => n1410);
   U5699 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxunsigned_output_9, Y
                           => n1429);
   U5700 : AOI22X1 port map( A0 => input_previous_1_10_port, A1 => n143, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_10_port, 
                           B1 => input_previous_1_17_port, Y => n4439);
   U5701 : XOR2X1 port map( A => n3694, B => input_previous_1_10_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_10_port);
   U5702 : NAND2X1 port map( A => n3679, B => n1293, Y => n3694);
   U5703 : AOI22X1 port map( A0 => input_previous_2_10_port, A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_10_port, 
                           B1 => input_previous_2_17_port, Y => n4492);
   U5704 : XOR2X1 port map( A => n3742, B => input_previous_2_10_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_10_port);
   U5705 : NAND2X1 port map( A => n3727, B => n1283, Y => n3742);
   U5706 : AOI22X1 port map( A0 => output_previous_2_10_port, A1 => n139, B0 =>
                           output_p2_times_a2_mul_componentxinput_A_inverted_10_port, 
                           B1 => output_previous_2_17_port, Y => n4598);
   U5707 : XOR2X1 port map( A => n3838, B => output_previous_2_10_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_10_port);
   U5708 : NAND2X1 port map( A => n3823, B => n1282, Y => n3838);
   U5709 : AOI22X1 port map( A0 => input_previous_0_10_port, A1 => n131, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_10_port, 
                           B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn88);
   U5710 : XOR2X1 port map( A => n3646, B => input_previous_0_10_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_10_port);
   U5711 : NAND2X1 port map( A => n3631, B => n1191, Y => n3646);
   U5712 : AOI22X1 port map( A0 => input_previous_1_11_port, A1 => n143, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_11_port, 
                           B1 => input_previous_1_17_port, Y => n4438);
   U5713 : XOR2X1 port map( A => n3692, B => input_previous_1_11_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_11_port);
   U5714 : AOI22X1 port map( A0 => input_previous_0_11_port, A1 => n131, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_11_port, 
                           B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn87);
   U5715 : XOR2X1 port map( A => n3644, B => input_previous_0_11_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_11_port);
   U5716 : NOR3X1 port map( A => input_previous_1_7_port, B => 
                           input_previous_1_8_port, C => n3681, Y => n3679);
   U5717 : NOR3X1 port map( A => input_previous_0_7_port, B => 
                           input_previous_0_8_port, C => n3633, Y => n3631);
   U5718 : NOR3X1 port map( A => input_previous_2_7_port, B => 
                           input_previous_2_8_port, C => n3729, Y => n3727);
   U5719 : NOR3X1 port map( A => output_previous_2_7_port, B => 
                           output_previous_2_8_port, C => n3825, Y => n3823);
   U5720 : NAND3BX1 port map( AN => input_previous_1_10_port, B => n1293, C => 
                           n3679, Y => n3692);
   U5721 : NAND3BX1 port map( AN => input_previous_0_10_port, B => n1191, C => 
                           n3631, Y => n3644);
   U5722 : OR3XL port map( A => input_previous_1_5_port, B => 
                           input_previous_1_6_port, C => n3683, Y => n3681);
   U5723 : OR3XL port map( A => input_previous_0_5_port, B => 
                           input_previous_0_6_port, C => n3635, Y => n3633);
   U5724 : OR3XL port map( A => input_previous_2_5_port, B => 
                           input_previous_2_6_port, C => n3731, Y => n3729);
   U5725 : OR3XL port map( A => output_previous_2_5_port, B => 
                           output_previous_2_6_port, C => n3827, Y => n3825);
   U5726 : OR3XL port map( A => input_previous_1_1_port, B => 
                           input_previous_1_2_port, C => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_0_port, Y 
                           => n3685);
   U5727 : OR3XL port map( A => input_previous_0_1_port, B => 
                           input_previous_0_2_port, C => 
                           input_times_b0_mul_componentxinput_A_inverted_0_port
                           , Y => n3637);
   U5728 : OR3XL port map( A => input_previous_2_1_port, B => 
                           input_previous_2_2_port, C => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_0_port, Y 
                           => n3733);
   U5729 : OR3XL port map( A => output_previous_2_1_port, B => 
                           output_previous_2_2_port, C => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_0_port, Y 
                           => n3829);
   U5730 : OR3XL port map( A => input_previous_1_3_port, B => 
                           input_previous_1_4_port, C => n3685, Y => n3683);
   U5731 : OR3XL port map( A => input_previous_0_3_port, B => 
                           input_previous_0_4_port, C => n3637, Y => n3635);
   U5732 : OR3XL port map( A => input_previous_2_3_port, B => 
                           input_previous_2_4_port, C => n3733, Y => n3731);
   U5733 : OR3XL port map( A => output_previous_2_3_port, B => 
                           output_previous_2_4_port, C => n3829, Y => n3827);
   U5734 : INVX1 port map( A => n4205, Y => n373);
   U5735 : AOI22X1 port map( A0 => n4203, A1 => 
                           input_p1_times_b1_div_componentxoutput_sign_gated_prev, 
                           B0 => n4204, B1 => n374, Y => n4205);
   U5736 : XNOR2X1 port map( A => n124, B => n333, Y => n4204);
   U5737 : INVX1 port map( A => n4261, Y => n375);
   U5738 : AOI22X1 port map( A0 => n4259, A1 => 
                           input_p2_times_b2_div_componentxoutput_sign_gated_prev, 
                           B0 => n4260, B1 => n376, Y => n4261);
   U5739 : XNOR2X1 port map( A => n128, B => n324, Y => n4260);
   U5740 : INVX1 port map( A => n4371, Y => n377);
   U5741 : AOI22X1 port map( A0 => n4369, A1 => 
                           output_p2_times_a2_div_componentxoutput_sign_gated_prev, 
                           B0 => n4370, B1 => n378, Y => n4371);
   U5742 : XNOR2X1 port map( A => n116, B => n351, Y => n4370);
   U5743 : INVX1 port map( A => input_times_b0_div_componentxn27, Y => n379);
   U5744 : AOI22X1 port map( A0 => input_times_b0_div_componentxn24, A1 => 
                           input_times_b0_div_componentxoutput_sign_gated_prev,
                           B0 => input_times_b0_div_componentxn25, B1 => n380, 
                           Y => input_times_b0_div_componentxn27);
   U5745 : XNOR2X1 port map( A => n120, B => n342, Y => 
                           input_times_b0_div_componentxn25);
   U5746 : BUFX3 port map( A => n4424, Y => n180);
   U5747 : AOI22X1 port map( A0 => input_previous_1_9_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_9_port, 
                           B1 => input_previous_1_17_port, Y => n4424);
   U5748 : XNOR2X1 port map( A => n3679, B => input_previous_1_9_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_9_port);
   U5749 : BUFX3 port map( A => n4477, Y => n201);
   U5750 : AOI22X1 port map( A0 => input_previous_2_9_port, A1 => n142, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_9_port, 
                           B1 => input_previous_2_17_port, Y => n4477);
   U5751 : XNOR2X1 port map( A => n3727, B => input_previous_2_9_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_9_port);
   U5752 : BUFX3 port map( A => n4583, Y => n243);
   U5753 : AOI22X1 port map( A0 => output_previous_2_9_port, A1 => n140, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_9_port, 
                           B1 => output_previous_2_17_port, Y => n4583);
   U5754 : XNOR2X1 port map( A => n3823, B => output_previous_2_9_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_9_port);
   U5755 : BUFX3 port map( A => input_times_b0_mul_componentxn73, Y => n271);
   U5756 : AOI22X1 port map( A0 => input_previous_0_9_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_9_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn73);
   U5757 : XNOR2X1 port map( A => n3631, B => input_previous_0_9_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_9_port
                           );
   U5758 : OAI2BB1X1 port map( A0N => 
                           input_p1_times_b1_div_componentxUDxshifted_substraction_result_0, 
                           A1N => n370, B0 => n1869, Y => n1889);
   U5759 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_16, 
                           A1 => n1870, B0 => 
                           input_p1_times_b1_div_componentxunsigned_A_17, B1 =>
                           n1871, Y => n1869);
   U5760 : NOR2BX1 port map( AN => 
                           input_p1_times_b1_div_componentxinput_A_inverted_17_port, B 
                           => n190, Y => 
                           input_p1_times_b1_div_componentxunsigned_A_17);
   U5761 : XOR2X1 port map( A => n3919, B => n123, Y => 
                           input_p1_times_b1_div_componentxinput_A_inverted_17_port);
   U5762 : OAI2BB1X1 port map( A0N => 
                           input_p2_times_b2_div_componentxUDxshifted_substraction_result_0, 
                           A1N => n369, B0 => n1979, Y => n1998);
   U5763 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_16, 
                           A1 => n1980, B0 => 
                           input_p2_times_b2_div_componentxunsigned_A_17, B1 =>
                           n1, Y => n1979);
   U5764 : NOR2BX1 port map( AN => 
                           input_p2_times_b2_div_componentxinput_A_inverted_17_port, B 
                           => n211, Y => 
                           input_p2_times_b2_div_componentxunsigned_A_17);
   U5765 : XOR2X1 port map( A => n3962, B => n127, Y => 
                           input_p2_times_b2_div_componentxinput_A_inverted_17_port);
   U5766 : OAI2BB1X1 port map( A0N => 
                           output_p2_times_a2_div_componentxUDxshifted_substraction_result_0, 
                           A1N => n368, B0 => n2198, Y => n2217);
   U5767 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_16, 
                           A1 => n2199, B0 => 
                           output_p2_times_a2_div_componentxunsigned_A_17, B1 
                           => n2090, Y => n2198);
   U5768 : NOR2BX1 port map( AN => 
                           output_p2_times_a2_div_componentxinput_A_inverted_17_port, B 
                           => n253, Y => 
                           output_p2_times_a2_div_componentxunsigned_A_17);
   U5769 : XOR2X1 port map( A => n4048, B => n115, Y => 
                           output_p2_times_a2_div_componentxinput_A_inverted_17_port);
   U5770 : OAI2BB1X1 port map( A0N => 
                           input_times_b0_div_componentxUDxshifted_substraction_result_0, 
                           A1N => n368, B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn2, 
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn22)
                           ;
   U5771 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_16, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => input_times_b0_div_componentxunsigned_A_17, B1
                           => n1871, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn2);
   U5772 : NOR2BX1 port map( AN => 
                           input_times_b0_div_componentxinput_A_inverted_17_port, B 
                           => n281, Y => 
                           input_times_b0_div_componentxunsigned_A_17);
   U5773 : XOR2X1 port map( A => n3876, B => n119, Y => 
                           input_times_b0_div_componentxinput_A_inverted_17_port);
   U5774 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_1, 
                           B0 => n1887, Y => n1905);
   U5775 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_0, 
                           A1 => n1870, B0 => n857, B1 => n1871, Y => n1887);
   U5776 : INVX1 port map( A => n4207, Y => n857);
   U5777 : AOI22X1 port map( A0 => n994, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_1_port, 
                           B1 => n124, Y => n4207);
   U5778 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_2, 
                           B0 => n1886, Y => n1904);
   U5779 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_1, 
                           A1 => n1870, B0 => n858, B1 => n1871, Y => n1886);
   U5780 : INVX1 port map( A => n4208, Y => n858);
   U5781 : AOI22X1 port map( A0 => n993, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_2_port, 
                           B1 => n124, Y => n4208);
   U5782 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_3, 
                           B0 => n1885, Y => n1903);
   U5783 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_2, 
                           A1 => n1870, B0 => n859, B1 => n1871, Y => n1885);
   U5784 : INVX1 port map( A => n4209, Y => n859);
   U5785 : AOI22X1 port map( A0 => n986, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_3_port, 
                           B1 => n124, Y => n4209);
   U5786 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_4, 
                           B0 => n1884, Y => n1902);
   U5787 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_3, 
                           A1 => n1870, B0 => n860, B1 => n1871, Y => n1884);
   U5788 : INVX1 port map( A => n4210, Y => n860);
   U5789 : AOI22X1 port map( A0 => n980, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_4_port, 
                           B1 => n124, Y => n4210);
   U5790 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_5, 
                           B0 => n1883, Y => n1901);
   U5791 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_4, 
                           A1 => n1870, B0 => n861, B1 => n1871, Y => n1883);
   U5792 : INVX1 port map( A => n4211, Y => n861);
   U5793 : AOI22X1 port map( A0 => n972, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_5_port, 
                           B1 => n124, Y => n4211);
   U5794 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_6, 
                           B0 => n1882, Y => n1900);
   U5795 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_5, 
                           A1 => n1870, B0 => n862, B1 => n1871, Y => n1882);
   U5796 : INVX1 port map( A => n4212, Y => n862);
   U5797 : AOI22X1 port map( A0 => n965, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_6_port, 
                           B1 => n124, Y => n4212);
   U5798 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_7, 
                           B0 => n1881, Y => n1899);
   U5799 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_6, 
                           A1 => n1870, B0 => n863, B1 => n1871, Y => n1881);
   U5800 : INVX1 port map( A => n4213, Y => n863);
   U5801 : AOI22X1 port map( A0 => n957, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_7_port, 
                           B1 => n124, Y => n4213);
   U5802 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_8, 
                           B0 => n1880, Y => n1898);
   U5803 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_7, 
                           A1 => n1870, B0 => n864, B1 => n1871, Y => n1880);
   U5804 : INVX1 port map( A => n4214, Y => n864);
   U5805 : AOI22X1 port map( A0 => n950, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_8_port, 
                           B1 => n124, Y => n4214);
   U5806 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_9, 
                           B0 => n1879, Y => n1897);
   U5807 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_8, 
                           A1 => n1870, B0 => n865, B1 => n1871, Y => n1879);
   U5808 : INVX1 port map( A => n4215, Y => n865);
   U5809 : AOI22X1 port map( A0 => n940, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_9_port, 
                           B1 => n123, Y => n4215);
   U5810 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_10, 
                           B0 => n1878, Y => n1896);
   U5811 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_9, 
                           A1 => n1870, B0 => n866, B1 => n1871, Y => n1878);
   U5812 : INVX1 port map( A => n4216, Y => n866);
   U5813 : AOI22X1 port map( A0 => n930, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_10_port, 
                           B1 => n123, Y => n4216);
   U5814 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_11, 
                           B0 => n1877, Y => n1895);
   U5815 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_10, 
                           A1 => n1870, B0 => n867, B1 => n1871, Y => n1877);
   U5816 : INVX1 port map( A => n4217, Y => n867);
   U5817 : AOI22X1 port map( A0 => n917, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_11_port, 
                           B1 => n123, Y => n4217);
   U5818 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_12, 
                           B0 => n1876, Y => n1894);
   U5819 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_11, 
                           A1 => n1870, B0 => n868, B1 => n1871, Y => n1876);
   U5820 : INVX1 port map( A => n4218, Y => n868);
   U5821 : AOI22X1 port map( A0 => n908, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_12_port, 
                           B1 => n123, Y => n4218);
   U5822 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_13, 
                           B0 => n1875, Y => n1893);
   U5823 : AOI22XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_12, 
                           A1 => n1870, B0 => n869, B1 => n1871, Y => n1875);
   U5824 : INVX1 port map( A => n4219, Y => n869);
   U5825 : AOI22X1 port map( A0 => n899, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_13_port, 
                           B1 => n123, Y => n4219);
   U5826 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_14, 
                           B0 => n1874, Y => n1892);
   U5827 : AOI22XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_13, 
                           A1 => n1870, B0 => n870, B1 => n1871, Y => n1874);
   U5828 : INVX1 port map( A => n4220, Y => n870);
   U5829 : AOI22X1 port map( A0 => n893, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_14_port, 
                           B1 => n123, Y => n4220);
   U5830 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_15, 
                           B0 => n1873, Y => n1891);
   U5831 : AOI22XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_14, 
                           A1 => n1870, B0 => n871, B1 => n1871, Y => n1873);
   U5832 : INVX1 port map( A => n4221, Y => n871);
   U5833 : AOI22X1 port map( A0 => n884, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_15_port, 
                           B1 => n123, Y => n4221);
   U5834 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_16, 
                           B0 => n1872, Y => n1890);
   U5835 : AOI22XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_15, 
                           A1 => n1870, B0 => n872, B1 => n1871, Y => n1872);
   U5836 : INVX1 port map( A => n4222, Y => n872);
   U5837 : AOI22X1 port map( A0 => n876, A1 => n190, B0 => 
                           input_p1_times_b1_div_componentxinput_A_inverted_16_port, 
                           B1 => n123, Y => n4222);
   U5838 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_1, 
                           B0 => n1996, Y => n2014);
   U5839 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_0, 
                           A1 => n1980, B0 => n1016, B1 => n1, Y => n1996);
   U5840 : INVX1 port map( A => n4263, Y => n1016);
   U5841 : AOI22X1 port map( A0 => n1153, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_1_port, 
                           B1 => n128, Y => n4263);
   U5842 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_2, 
                           B0 => n1995, Y => n2013);
   U5843 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_1, 
                           A1 => n1980, B0 => n1017, B1 => n1, Y => n1995);
   U5844 : INVX1 port map( A => n4264, Y => n1017);
   U5845 : AOI22X1 port map( A0 => n1152, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_2_port, 
                           B1 => n128, Y => n4264);
   U5846 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_3, 
                           B0 => n1994, Y => n2012);
   U5847 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_2, 
                           A1 => n1980, B0 => n1018, B1 => n1, Y => n1994);
   U5848 : INVX1 port map( A => n4265, Y => n1018);
   U5849 : AOI22X1 port map( A0 => n1145, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_3_port, 
                           B1 => n128, Y => n4265);
   U5850 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_4, 
                           B0 => n1993, Y => n2011);
   U5851 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_3, 
                           A1 => n1980, B0 => n1019, B1 => n1, Y => n1993);
   U5852 : INVX1 port map( A => n4266, Y => n1019);
   U5853 : AOI22X1 port map( A0 => n1139, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_4_port, 
                           B1 => n128, Y => n4266);
   U5854 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_5, 
                           B0 => n1992, Y => n2010);
   U5855 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_4, 
                           A1 => n1980, B0 => n1020, B1 => n1, Y => n1992);
   U5856 : INVX1 port map( A => n4267, Y => n1020);
   U5857 : AOI22X1 port map( A0 => n1131, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_5_port, 
                           B1 => n128, Y => n4267);
   U5858 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_6, 
                           B0 => n1991, Y => n2009);
   U5859 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_5, 
                           A1 => n1980, B0 => n1021, B1 => n1, Y => n1991);
   U5860 : INVX1 port map( A => n4268, Y => n1021);
   U5861 : AOI22X1 port map( A0 => n1124, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_6_port, 
                           B1 => n128, Y => n4268);
   U5862 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_7, 
                           B0 => n1990, Y => n2008);
   U5863 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_6, 
                           A1 => n1980, B0 => n1022, B1 => n1, Y => n1990);
   U5864 : INVX1 port map( A => n4269, Y => n1022);
   U5865 : AOI22X1 port map( A0 => n1116, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_7_port, 
                           B1 => n128, Y => n4269);
   U5866 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_8, 
                           B0 => n1989, Y => n2007);
   U5867 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_7, 
                           A1 => n1980, B0 => n1023, B1 => n1, Y => n1989);
   U5868 : INVX1 port map( A => n4270, Y => n1023);
   U5869 : AOI22X1 port map( A0 => n1109, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_8_port, 
                           B1 => n128, Y => n4270);
   U5870 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_9, 
                           B0 => n1988, Y => n2006);
   U5871 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_8, 
                           A1 => n1980, B0 => n1024, B1 => n1, Y => n1988);
   U5872 : INVX1 port map( A => n4271, Y => n1024);
   U5873 : AOI22X1 port map( A0 => n1099, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_9_port, 
                           B1 => n127, Y => n4271);
   U5874 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_10, 
                           B0 => n1987, Y => n2005);
   U5875 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_9, 
                           A1 => n1980, B0 => n1025, B1 => n1, Y => n1987);
   U5876 : INVX1 port map( A => n4272, Y => n1025);
   U5877 : AOI22X1 port map( A0 => n1089, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_10_port, 
                           B1 => n127, Y => n4272);
   U5878 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_11, 
                           B0 => n1986, Y => n2004);
   U5879 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_10, 
                           A1 => n1980, B0 => n1026, B1 => n1, Y => n1986);
   U5880 : INVX1 port map( A => n4273, Y => n1026);
   U5881 : AOI22X1 port map( A0 => n1076, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_11_port, 
                           B1 => n127, Y => n4273);
   U5882 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_12, 
                           B0 => n1985, Y => n2003);
   U5883 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_11, 
                           A1 => n1980, B0 => n1027, B1 => n1, Y => n1985);
   U5884 : INVX1 port map( A => n4274, Y => n1027);
   U5885 : AOI22X1 port map( A0 => n1067, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_12_port, 
                           B1 => n127, Y => n4274);
   U5886 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_13, 
                           B0 => n1984, Y => n2002);
   U5887 : AOI22XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_12, 
                           A1 => n1980, B0 => n1028, B1 => n1, Y => n1984);
   U5888 : INVX1 port map( A => n4275, Y => n1028);
   U5889 : AOI22X1 port map( A0 => n1058, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_13_port, 
                           B1 => n127, Y => n4275);
   U5890 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_14, 
                           B0 => n1983, Y => n2001);
   U5891 : AOI22XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_13, 
                           A1 => n1980, B0 => n1029, B1 => n1, Y => n1983);
   U5892 : INVX1 port map( A => n4276, Y => n1029);
   U5893 : AOI22X1 port map( A0 => n1052, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_14_port, 
                           B1 => n127, Y => n4276);
   U5894 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_15, 
                           B0 => n1982, Y => n2000);
   U5895 : AOI22XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_14, 
                           A1 => n1980, B0 => n1030, B1 => n1, Y => n1982);
   U5896 : INVX1 port map( A => n4277, Y => n1030);
   U5897 : AOI22X1 port map( A0 => n1043, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_15_port, 
                           B1 => n127, Y => n4277);
   U5898 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_16, 
                           B0 => n1981, Y => n1999);
   U5899 : AOI22XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_15, 
                           A1 => n1980, B0 => n1031, B1 => n1, Y => n1981);
   U5900 : INVX1 port map( A => n4278, Y => n1031);
   U5901 : AOI22X1 port map( A0 => n1035, A1 => n211, B0 => 
                           input_p2_times_b2_div_componentxinput_A_inverted_16_port, 
                           B1 => n127, Y => n4278);
   U5902 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_1, 
                           B0 => n2215, Y => n2233);
   U5903 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_0, 
                           A1 => n2199, B0 => n539, B1 => n1871, Y => n2215);
   U5904 : INVX1 port map( A => n4373, Y => n539);
   U5905 : AOI22X1 port map( A0 => n676, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_1_port, 
                           B1 => n116, Y => n4373);
   U5906 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_2, 
                           B0 => n2214, Y => n2232);
   U5907 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_1, 
                           A1 => n2199, B0 => n540, B1 => n1, Y => n2214);
   U5908 : INVX1 port map( A => n4374, Y => n540);
   U5909 : AOI22X1 port map( A0 => n675, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_2_port, 
                           B1 => n116, Y => n4374);
   U5910 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_3, 
                           B0 => n2213, Y => n2231);
   U5911 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_2, 
                           A1 => n2199, B0 => n541, B1 => n2090, Y => n2213);
   U5912 : INVX1 port map( A => n4375, Y => n541);
   U5913 : AOI22X1 port map( A0 => n668, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_3_port, 
                           B1 => n116, Y => n4375);
   U5914 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_4, 
                           B0 => n2212, Y => n2230);
   U5915 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_3, 
                           A1 => n2199, B0 => n542, B1 => n1871, Y => n2212);
   U5916 : INVX1 port map( A => n4376, Y => n542);
   U5917 : AOI22X1 port map( A0 => n662, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_4_port, 
                           B1 => n116, Y => n4376);
   U5918 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_5, 
                           B0 => n2211, Y => n2229);
   U5919 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_4, 
                           A1 => n2199, B0 => n543, B1 => n1, Y => n2211);
   U5920 : INVX1 port map( A => n4377, Y => n543);
   U5921 : AOI22X1 port map( A0 => n654, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_5_port, 
                           B1 => n116, Y => n4377);
   U5922 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_6, 
                           B0 => n2210, Y => n2228);
   U5923 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_5, 
                           A1 => n2199, B0 => n544, B1 => n2090, Y => n2210);
   U5924 : INVX1 port map( A => n4378, Y => n544);
   U5925 : AOI22X1 port map( A0 => n647, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_6_port, 
                           B1 => n116, Y => n4378);
   U5926 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_7, 
                           B0 => n2209, Y => n2227);
   U5927 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_6, 
                           A1 => n2199, B0 => n545, B1 => n1871, Y => n2209);
   U5928 : INVX1 port map( A => n4379, Y => n545);
   U5929 : AOI22X1 port map( A0 => n639, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_7_port, 
                           B1 => n116, Y => n4379);
   U5930 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_8, 
                           B0 => n2208, Y => n2226);
   U5931 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_7, 
                           A1 => n2199, B0 => n546, B1 => n1, Y => n2208);
   U5932 : INVX1 port map( A => n4380, Y => n546);
   U5933 : AOI22X1 port map( A0 => n632, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_8_port, 
                           B1 => n116, Y => n4380);
   U5934 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_9, 
                           B0 => n2207, Y => n2225);
   U5935 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_8, 
                           A1 => n2199, B0 => n547, B1 => n2090, Y => n2207);
   U5936 : INVX1 port map( A => n4381, Y => n547);
   U5937 : AOI22X1 port map( A0 => n622, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_9_port, 
                           B1 => n115, Y => n4381);
   U5938 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_10, 
                           B0 => n2206, Y => n2224);
   U5939 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_9, 
                           A1 => n2199, B0 => n548, B1 => n1871, Y => n2206);
   U5940 : INVX1 port map( A => n4382, Y => n548);
   U5941 : AOI22X1 port map( A0 => n612, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_10_port, 
                           B1 => n115, Y => n4382);
   U5942 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_11, 
                           B0 => n2205, Y => n2223);
   U5943 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_10, 
                           A1 => n2199, B0 => n549, B1 => n1, Y => n2205);
   U5944 : INVX1 port map( A => n4383, Y => n549);
   U5945 : AOI22X1 port map( A0 => n599, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_11_port, 
                           B1 => n115, Y => n4383);
   U5946 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_12, 
                           B0 => n2204, Y => n2222);
   U5947 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_11, 
                           A1 => n2199, B0 => n550, B1 => n2090, Y => n2204);
   U5948 : INVX1 port map( A => n4384, Y => n550);
   U5949 : AOI22X1 port map( A0 => n590, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_12_port, 
                           B1 => n115, Y => n4384);
   U5950 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_13, 
                           B0 => n2203, Y => n2221);
   U5951 : AOI22XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_12, 
                           A1 => n2199, B0 => n551, B1 => n1, Y => n2203);
   U5952 : INVX1 port map( A => n4385, Y => n551);
   U5953 : AOI22X1 port map( A0 => n581, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_13_port, 
                           B1 => n115, Y => n4385);
   U5954 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_14, 
                           B0 => n2202, Y => n2220);
   U5955 : AOI22XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_13, 
                           A1 => n2199, B0 => n552, B1 => n2090, Y => n2202);
   U5956 : INVX1 port map( A => n4386, Y => n552);
   U5957 : AOI22X1 port map( A0 => n575, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_14_port, 
                           B1 => n115, Y => n4386);
   U5958 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_15, 
                           B0 => n2201, Y => n2219);
   U5959 : AOI22XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_14, 
                           A1 => n2199, B0 => n553, B1 => n1871, Y => n2201);
   U5960 : INVX1 port map( A => n4387, Y => n553);
   U5961 : AOI22X1 port map( A0 => n566, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_15_port, 
                           B1 => n115, Y => n4387);
   U5962 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_16, 
                           B0 => n2200, Y => n2218);
   U5963 : AOI22XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_15, 
                           A1 => n2199, B0 => n554, B1 => n1, Y => n2200);
   U5964 : INVX1 port map( A => n4388, Y => n554);
   U5965 : AOI22X1 port map( A0 => n558, A1 => n253, B0 => 
                           output_p2_times_a2_div_componentxinput_A_inverted_16_port, 
                           B1 => n115, Y => n4388);
   U5966 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_1, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn20,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn38)
                           ;
   U5967 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_0, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n698, B1 => n1, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn20)
                           ;
   U5968 : INVX1 port map( A => input_times_b0_div_componentxn29, Y => n698);
   U5969 : AOI22X1 port map( A0 => n835, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_1_port
                           , B1 => n120, Y => input_times_b0_div_componentxn29)
                           ;
   U5970 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_2, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn19,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn37)
                           ;
   U5971 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_1, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n699, B1 => n2090, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn19)
                           ;
   U5972 : INVX1 port map( A => input_times_b0_div_componentxn30, Y => n699);
   U5973 : AOI22X1 port map( A0 => n834, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_2_port
                           , B1 => n120, Y => input_times_b0_div_componentxn30)
                           ;
   U5974 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_3, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn18,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn36)
                           ;
   U5975 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_2, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n700, B1 => n2090, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn18)
                           ;
   U5976 : INVX1 port map( A => input_times_b0_div_componentxn31, Y => n700);
   U5977 : AOI22X1 port map( A0 => n827, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_3_port
                           , B1 => n120, Y => input_times_b0_div_componentxn31)
                           ;
   U5978 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_4, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn17,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn35)
                           ;
   U5979 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_3, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n701, B1 => n1871, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn17)
                           ;
   U5980 : INVX1 port map( A => input_times_b0_div_componentxn32, Y => n701);
   U5981 : AOI22X1 port map( A0 => n821, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_4_port
                           , B1 => n120, Y => input_times_b0_div_componentxn32)
                           ;
   U5982 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_5, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn16,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn34)
                           ;
   U5983 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_4, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n702, B1 => n1, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn16)
                           ;
   U5984 : INVX1 port map( A => input_times_b0_div_componentxn33, Y => n702);
   U5985 : AOI22X1 port map( A0 => n813, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_5_port
                           , B1 => n120, Y => input_times_b0_div_componentxn33)
                           ;
   U5986 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_6, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn15,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn33)
                           ;
   U5987 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_5, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n703, B1 => n2090, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn15)
                           ;
   U5988 : INVX1 port map( A => input_times_b0_div_componentxn34, Y => n703);
   U5989 : AOI22X1 port map( A0 => n806, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_6_port
                           , B1 => n120, Y => input_times_b0_div_componentxn34)
                           ;
   U5990 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_7, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn14,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn32)
                           ;
   U5991 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_6, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n704, B1 => n1871, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn14)
                           ;
   U5992 : INVX1 port map( A => input_times_b0_div_componentxn35, Y => n704);
   U5993 : AOI22X1 port map( A0 => n798, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_7_port
                           , B1 => n120, Y => input_times_b0_div_componentxn35)
                           ;
   U5994 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_8, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn13,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn31)
                           ;
   U5995 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_7, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n705, B1 => n1871, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn13)
                           ;
   U5996 : INVX1 port map( A => input_times_b0_div_componentxn36, Y => n705);
   U5997 : AOI22X1 port map( A0 => n791, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_8_port
                           , B1 => n120, Y => input_times_b0_div_componentxn36)
                           ;
   U5998 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_9, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn12,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn30)
                           ;
   U5999 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_8, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n706, B1 => n1, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn12)
                           ;
   U6000 : INVX1 port map( A => input_times_b0_div_componentxn37, Y => n706);
   U6001 : AOI22X1 port map( A0 => n781, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_9_port
                           , B1 => n119, Y => input_times_b0_div_componentxn37)
                           ;
   U6002 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_10, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn11,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn29)
                           ;
   U6003 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_9, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n707, B1 => n2090, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn11)
                           ;
   U6004 : INVX1 port map( A => input_times_b0_div_componentxn38, Y => n707);
   U6005 : AOI22X1 port map( A0 => n771, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_10_port, 
                           B1 => n119, Y => input_times_b0_div_componentxn38);
   U6006 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_11, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn10,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn28)
                           ;
   U6007 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_10, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n708, B1 => n1, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn10)
                           ;
   U6008 : INVX1 port map( A => input_times_b0_div_componentxn39, Y => n708);
   U6009 : AOI22X1 port map( A0 => n758, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_11_port, 
                           B1 => n119, Y => input_times_b0_div_componentxn39);
   U6010 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_12, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn9, 
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn27)
                           ;
   U6011 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_11, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n709, B1 => n1871, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn9);
   U6012 : INVX1 port map( A => input_times_b0_div_componentxn40, Y => n709);
   U6013 : AOI22X1 port map( A0 => n749, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_12_port, 
                           B1 => n119, Y => input_times_b0_div_componentxn40);
   U6014 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_13, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn8, 
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn26)
                           ;
   U6015 : AOI22XL port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_12, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n710, B1 => n1871, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn8);
   U6016 : INVX1 port map( A => input_times_b0_div_componentxn41, Y => n710);
   U6017 : AOI22X1 port map( A0 => n740, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_13_port, 
                           B1 => n119, Y => input_times_b0_div_componentxn41);
   U6018 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_14, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn7, 
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn25)
                           ;
   U6019 : AOI22XL port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_13, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n711, B1 => n1, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn7);
   U6020 : INVX1 port map( A => input_times_b0_div_componentxn42, Y => n711);
   U6021 : AOI22X1 port map( A0 => n734, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_14_port, 
                           B1 => n119, Y => input_times_b0_div_componentxn42);
   U6022 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_15, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn6, 
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn24)
                           ;
   U6023 : AOI22XL port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_14, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n712, B1 => n2090, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn6);
   U6024 : INVX1 port map( A => input_times_b0_div_componentxn43, Y => n712);
   U6025 : AOI22X1 port map( A0 => n725, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_15_port, 
                           B1 => n119, Y => input_times_b0_div_componentxn43);
   U6026 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_16, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn5, 
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn23)
                           ;
   U6027 : AOI22XL port map( A0 => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_15, 
                           A1 => 
                           input_times_b0_div_componentxUDxinput_containerxn3, 
                           B0 => n713, B1 => n2090, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn5);
   U6028 : INVX1 port map( A => input_times_b0_div_componentxn44, Y => n713);
   U6029 : AOI22X1 port map( A0 => n717, A1 => n281, B0 => 
                           input_times_b0_div_componentxinput_A_inverted_16_port, 
                           B1 => n119, Y => input_times_b0_div_componentxn44);
   U6030 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxinput_containerxparallel_out_0, 
                           B0 => n1888, Y => n1906);
   U6031 : NAND2XL port map( A => n856, B => n1871, Y => n1888);
   U6032 : INVX1 port map( A => n4206, Y => n856);
   U6033 : AOI22X1 port map( A0 => n995, A1 => n190, B0 => n995, B1 => n124, Y 
                           => n4206);
   U6034 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxinput_containerxparallel_out_0, 
                           B0 => n1997, Y => n2015);
   U6035 : NAND2XL port map( A => n1015, B => n1, Y => n1997);
   U6036 : INVX1 port map( A => n4262, Y => n1015);
   U6037 : AOI22X1 port map( A0 => n1154, A1 => n211, B0 => n1154, B1 => n128, 
                           Y => n4262);
   U6038 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p2_times_a2_div_componentxUDxinput_containerxparallel_out_0, 
                           B0 => n2216, Y => n2234);
   U6039 : NAND2XL port map( A => n538, B => n1871, Y => n2216);
   U6040 : INVX1 port map( A => n4372, Y => n538);
   U6041 : AOI22X1 port map( A0 => n677, A1 => n253, B0 => n677, B1 => n116, Y 
                           => n4372);
   U6042 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_times_b0_div_componentxUDxinput_containerxparallel_out_0, 
                           B0 => 
                           input_times_b0_div_componentxUDxinput_containerxn21,
                           Y => 
                           input_times_b0_div_componentxUDxinput_containerxn40)
                           ;
   U6043 : NAND2XL port map( A => n697, B => n1, Y => 
                           input_times_b0_div_componentxUDxinput_containerxn21)
                           ;
   U6044 : INVX1 port map( A => input_times_b0_div_componentxn28, Y => n697);
   U6045 : AOI22X1 port map( A0 => n836, A1 => n281, B0 => n836, B1 => n120, Y 
                           => input_times_b0_div_componentxn28);
   U6046 : AOI22X1 port map( A0 => input_previous_2_11_port, A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_11_port, 
                           B1 => input_previous_2_17_port, Y => n4491);
   U6047 : XOR2X1 port map( A => n3740, B => input_previous_2_11_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_11_port);
   U6048 : AOI22X1 port map( A0 => output_previous_2_11_port, A1 => n139, B0 =>
                           output_p2_times_a2_mul_componentxinput_A_inverted_11_port, 
                           B1 => output_previous_2_17_port, Y => n4597);
   U6049 : XOR2X1 port map( A => n3836, B => output_previous_2_11_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_11_port);
   U6050 : AOI22X1 port map( A0 => input_previous_2_12_port, A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_12_port, 
                           B1 => input_previous_2_17_port, Y => n4490);
   U6051 : XOR2X1 port map( A => n3741, B => input_previous_2_12_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_12_port);
   U6052 : OR2X2 port map( A => n3740, B => input_previous_2_11_port, Y => 
                           n3741);
   U6053 : AOI22X1 port map( A0 => output_previous_2_12_port, A1 => n139, B0 =>
                           output_p2_times_a2_mul_componentxinput_A_inverted_12_port, 
                           B1 => output_previous_2_17_port, Y => n4596);
   U6054 : XOR2X1 port map( A => n3837, B => output_previous_2_12_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_12_port);
   U6055 : OR2X2 port map( A => n3836, B => output_previous_2_11_port, Y => 
                           n3837);
   U6056 : AOI22X1 port map( A0 => input_previous_1_13_port, A1 => n143, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_13_port, 
                           B1 => input_previous_1_17_port, Y => n4436);
   U6057 : XOR2X1 port map( A => n3690, B => input_previous_1_13_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_13_port);
   U6058 : AOI22X1 port map( A0 => input_previous_2_13_port, A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_13_port, 
                           B1 => input_previous_2_17_port, Y => n4489);
   U6059 : XOR2X1 port map( A => n3738, B => input_previous_2_13_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_13_port);
   U6060 : AOI22X1 port map( A0 => output_previous_2_13_port, A1 => n139, B0 =>
                           output_p2_times_a2_mul_componentxinput_A_inverted_13_port, 
                           B1 => output_previous_2_17_port, Y => n4595);
   U6061 : XOR2X1 port map( A => n3834, B => output_previous_2_13_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_13_port);
   U6062 : AOI22X1 port map( A0 => input_previous_0_13_port, A1 => n131, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_13_port, 
                           B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn85);
   U6063 : XOR2X1 port map( A => n3642, B => input_previous_0_13_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_13_port);
   U6064 : AOI22X1 port map( A0 => input_previous_1_14_port, A1 => n143, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_14_port, 
                           B1 => input_previous_1_17_port, Y => n4435);
   U6065 : XOR2X1 port map( A => n3691, B => input_previous_1_14_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_14_port);
   U6066 : OR2X2 port map( A => input_previous_1_13_port, B => n3690, Y => 
                           n3691);
   U6067 : AOI22X1 port map( A0 => input_previous_2_14_port, A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_14_port, 
                           B1 => input_previous_2_17_port, Y => n4488);
   U6068 : XOR2X1 port map( A => n3739, B => input_previous_2_14_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_14_port);
   U6069 : OR2X2 port map( A => input_previous_2_13_port, B => n3738, Y => 
                           n3739);
   U6070 : AOI22X1 port map( A0 => output_previous_2_14_port, A1 => n139, B0 =>
                           output_p2_times_a2_mul_componentxinput_A_inverted_14_port, 
                           B1 => output_previous_2_17_port, Y => n4594);
   U6071 : XOR2X1 port map( A => n3835, B => output_previous_2_14_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_14_port);
   U6072 : OR2X2 port map( A => output_previous_2_13_port, B => n3834, Y => 
                           n3835);
   U6073 : AOI22X1 port map( A0 => input_previous_0_14_port, A1 => n131, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_14_port, 
                           B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn84);
   U6074 : XOR2X1 port map( A => n3643, B => input_previous_0_14_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_14_port);
   U6075 : OR2X2 port map( A => input_previous_0_13_port, B => n3642, Y => 
                           n3643);
   U6076 : AOI22X1 port map( A0 => input_previous_2_15_port, A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_15_port, 
                           B1 => input_previous_2_17_port, Y => n4487);
   U6077 : XNOR2X1 port map( A => n3737, B => input_previous_2_15_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_15_port);
   U6078 : AOI22X1 port map( A0 => output_previous_2_15_port, A1 => n139, B0 =>
                           output_p2_times_a2_mul_componentxinput_A_inverted_15_port, 
                           B1 => output_previous_2_17_port, Y => n4593);
   U6079 : XNOR2X1 port map( A => n3833, B => output_previous_2_15_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_15_port);
   U6080 : NOR3X1 port map( A => input_previous_1_13_port, B => 
                           input_previous_1_14_port, C => n3690, Y => n3689);
   U6081 : NOR3X1 port map( A => input_previous_0_13_port, B => 
                           input_previous_0_14_port, C => n3642, Y => n3641);
   U6082 : NOR3X1 port map( A => input_previous_2_13_port, B => 
                           input_previous_2_14_port, C => n3738, Y => n3737);
   U6083 : NOR3X1 port map( A => output_previous_2_13_port, B => 
                           output_previous_2_14_port, C => n3834, Y => n3833);
   U6084 : BUFX3 port map( A => n4429, Y => n185);
   U6085 : AOI22X1 port map( A0 => input_previous_1_4_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_4_port, 
                           B1 => input_previous_1_17_port, Y => n4429);
   U6086 : XOR2X1 port map( A => n3684, B => input_previous_1_4_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_4_port);
   U6087 : OR2X2 port map( A => input_previous_1_3_port, B => n3685, Y => n3684
                           );
   U6088 : BUFX3 port map( A => input_times_b0_mul_componentxn78, Y => n276);
   U6089 : AOI22X1 port map( A0 => input_previous_0_4_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_4_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn78);
   U6090 : XOR2X1 port map( A => n3636, B => input_previous_0_4_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_4_port
                           );
   U6091 : OR2X2 port map( A => input_previous_0_3_port, B => n3637, Y => n3636
                           );
   U6092 : NAND3BX1 port map( AN => input_previous_2_10_port, B => n1283, C => 
                           n3727, Y => n3740);
   U6093 : NAND3BX1 port map( AN => output_previous_2_10_port, B => n1282, C =>
                           n3823, Y => n3836);
   U6094 : OR3XL port map( A => input_previous_1_11_port, B => 
                           input_previous_1_12_port, C => n3692, Y => n3690);
   U6095 : OR3XL port map( A => input_previous_0_11_port, B => 
                           input_previous_0_12_port, C => n3644, Y => n3642);
   U6096 : OR3XL port map( A => input_previous_2_11_port, B => 
                           input_previous_2_12_port, C => n3740, Y => n3738);
   U6097 : OR3XL port map( A => output_previous_2_11_port, B => 
                           output_previous_2_12_port, C => n3836, Y => n3834);
   U6098 : BUFX3 port map( A => n4440, Y => n189);
   U6099 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_0_port, 
                           A1 => n143, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_0_port, 
                           B1 => input_previous_1_17_port, Y => n4440);
   U6100 : BUFX3 port map( A => n4493, Y => n210);
   U6101 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_0_port, 
                           A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_0_port, 
                           B1 => input_previous_2_17_port, Y => n4493);
   U6102 : BUFX3 port map( A => n4599, Y => n252);
   U6103 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_0_port, 
                           A1 => n139, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_0_port, 
                           B1 => output_previous_2_17_port, Y => n4599);
   U6104 : BUFX3 port map( A => input_times_b0_mul_componentxn89, Y => n280);
   U6105 : AOI22X1 port map( A0 => 
                           input_times_b0_mul_componentxinput_A_inverted_0_port
                           , A1 => n131, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_0_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn89);
   U6106 : BUFX3 port map( A => n4432, Y => n188);
   U6107 : AOI22X1 port map( A0 => input_previous_1_1_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_1_port, 
                           B1 => input_previous_1_17_port, Y => n4432);
   U6108 : XOR2X1 port map( A => input_previous_1_1_port, B => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_0_port, Y 
                           => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_1_port);
   U6109 : BUFX3 port map( A => n4485, Y => n209);
   U6110 : AOI22X1 port map( A0 => input_previous_2_1_port, A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_1_port, 
                           B1 => input_previous_2_17_port, Y => n4485);
   U6111 : XOR2X1 port map( A => input_previous_2_1_port, B => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_0_port, Y 
                           => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_1_port);
   U6112 : BUFX3 port map( A => n4591, Y => n251);
   U6113 : AOI22X1 port map( A0 => output_previous_2_1_port, A1 => n139, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_1_port, 
                           B1 => output_previous_2_17_port, Y => n4591);
   U6114 : XOR2X1 port map( A => output_previous_2_1_port, B => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_0_port, Y 
                           => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_1_port);
   U6115 : BUFX3 port map( A => input_times_b0_mul_componentxn81, Y => n279);
   U6116 : AOI22X1 port map( A0 => input_previous_0_1_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_1_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn81);
   U6117 : XOR2X1 port map( A => input_previous_0_1_port, B => 
                           input_times_b0_mul_componentxinput_A_inverted_0_port
                           , Y => 
                           input_times_b0_mul_componentxinput_A_inverted_1_port
                           );
   U6118 : BUFX3 port map( A => n4431, Y => n187);
   U6119 : AOI22X1 port map( A0 => input_previous_1_2_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_2_port, 
                           B1 => input_previous_1_17_port, Y => n4431);
   U6120 : XNOR2X1 port map( A => input_previous_1_2_port, B => n3686, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_2_port);
   U6121 : NOR2X1 port map( A => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_0_port, B 
                           => input_previous_1_1_port, Y => n3686);
   U6122 : BUFX3 port map( A => n4484, Y => n208);
   U6123 : AOI22X1 port map( A0 => input_previous_2_2_port, A1 => n142, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_2_port, 
                           B1 => input_previous_2_17_port, Y => n4484);
   U6124 : XNOR2X1 port map( A => input_previous_2_2_port, B => n3734, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_2_port);
   U6125 : NOR2X1 port map( A => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_0_port, B 
                           => input_previous_2_1_port, Y => n3734);
   U6126 : BUFX3 port map( A => n4590, Y => n250);
   U6127 : AOI22X1 port map( A0 => output_previous_2_2_port, A1 => n140, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_2_port, 
                           B1 => output_previous_2_17_port, Y => n4590);
   U6128 : XNOR2X1 port map( A => output_previous_2_2_port, B => n3830, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_2_port);
   U6129 : NOR2X1 port map( A => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_0_port, B 
                           => output_previous_2_1_port, Y => n3830);
   U6130 : BUFX3 port map( A => input_times_b0_mul_componentxn80, Y => n278);
   U6131 : AOI22X1 port map( A0 => input_previous_0_2_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_2_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn80);
   U6132 : XNOR2X1 port map( A => input_previous_0_2_port, B => n3638, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_2_port
                           );
   U6133 : NOR2X1 port map( A => 
                           input_times_b0_mul_componentxinput_A_inverted_0_port
                           , B => input_previous_0_1_port, Y => n3638);
   U6134 : BUFX3 port map( A => n4430, Y => n186);
   U6135 : AOI22X1 port map( A0 => input_previous_1_3_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_3_port, 
                           B1 => input_previous_1_17_port, Y => n4430);
   U6136 : XOR2X1 port map( A => n3685, B => input_previous_1_3_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_3_port);
   U6137 : BUFX3 port map( A => input_times_b0_mul_componentxn79, Y => n277);
   U6138 : AOI22X1 port map( A0 => input_previous_0_3_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_3_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn79);
   U6139 : XOR2X1 port map( A => n3637, B => input_previous_0_3_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_3_port
                           );
   U6140 : BUFX3 port map( A => n4428, Y => n184);
   U6141 : AOI22X1 port map( A0 => input_previous_1_5_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_5_port, 
                           B1 => input_previous_1_17_port, Y => n4428);
   U6142 : XOR2X1 port map( A => n3683, B => input_previous_1_5_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_5_port);
   U6143 : BUFX3 port map( A => n4481, Y => n205);
   U6144 : AOI22X1 port map( A0 => input_previous_2_5_port, A1 => n142, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_5_port, 
                           B1 => input_previous_2_17_port, Y => n4481);
   U6145 : XOR2X1 port map( A => n3731, B => input_previous_2_5_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_5_port);
   U6146 : BUFX3 port map( A => n4587, Y => n247);
   U6147 : AOI22X1 port map( A0 => output_previous_2_5_port, A1 => n140, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_5_port, 
                           B1 => output_previous_2_17_port, Y => n4587);
   U6148 : XOR2X1 port map( A => n3827, B => output_previous_2_5_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_5_port);
   U6149 : BUFX3 port map( A => input_times_b0_mul_componentxn77, Y => n275);
   U6150 : AOI22X1 port map( A0 => input_previous_0_5_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_5_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn77);
   U6151 : XOR2X1 port map( A => n3635, B => input_previous_0_5_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_5_port
                           );
   U6152 : BUFX3 port map( A => n4427, Y => n183);
   U6153 : AOI22X1 port map( A0 => input_previous_1_6_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_6_port, 
                           B1 => input_previous_1_17_port, Y => n4427);
   U6154 : XOR2X1 port map( A => n3682, B => input_previous_1_6_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_6_port);
   U6155 : OR2X2 port map( A => input_previous_1_5_port, B => n3683, Y => n3682
                           );
   U6156 : BUFX3 port map( A => n4480, Y => n204);
   U6157 : AOI22X1 port map( A0 => input_previous_2_6_port, A1 => n142, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_6_port, 
                           B1 => input_previous_2_17_port, Y => n4480);
   U6158 : XOR2X1 port map( A => n3730, B => input_previous_2_6_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_6_port);
   U6159 : OR2X2 port map( A => input_previous_2_5_port, B => n3731, Y => n3730
                           );
   U6160 : BUFX3 port map( A => n4586, Y => n246);
   U6161 : AOI22X1 port map( A0 => output_previous_2_6_port, A1 => n140, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_6_port, 
                           B1 => output_previous_2_17_port, Y => n4586);
   U6162 : XOR2X1 port map( A => n3826, B => output_previous_2_6_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_6_port);
   U6163 : OR2X2 port map( A => output_previous_2_5_port, B => n3827, Y => 
                           n3826);
   U6164 : BUFX3 port map( A => input_times_b0_mul_componentxn76, Y => n274);
   U6165 : AOI22X1 port map( A0 => input_previous_0_6_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_6_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn76);
   U6166 : XOR2X1 port map( A => n3634, B => input_previous_0_6_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_6_port
                           );
   U6167 : OR2X2 port map( A => input_previous_0_5_port, B => n3635, Y => n3634
                           );
   U6168 : BUFX3 port map( A => n4426, Y => n182);
   U6169 : AOI22X1 port map( A0 => input_previous_1_7_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_7_port, 
                           B1 => input_previous_1_17_port, Y => n4426);
   U6170 : XOR2X1 port map( A => n3681, B => input_previous_1_7_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_7_port);
   U6171 : BUFX3 port map( A => n4479, Y => n203);
   U6172 : AOI22X1 port map( A0 => input_previous_2_7_port, A1 => n142, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_7_port, 
                           B1 => input_previous_2_17_port, Y => n4479);
   U6173 : XOR2X1 port map( A => n3729, B => input_previous_2_7_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_7_port);
   U6174 : BUFX3 port map( A => n4585, Y => n245);
   U6175 : AOI22X1 port map( A0 => output_previous_2_7_port, A1 => n140, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_7_port, 
                           B1 => output_previous_2_17_port, Y => n4585);
   U6176 : XOR2X1 port map( A => n3825, B => output_previous_2_7_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_7_port);
   U6177 : BUFX3 port map( A => input_times_b0_mul_componentxn75, Y => n273);
   U6178 : AOI22X1 port map( A0 => input_previous_0_7_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_7_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn75);
   U6179 : XOR2X1 port map( A => n3633, B => input_previous_0_7_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_7_port
                           );
   U6180 : AOI22X1 port map( A0 => input_previous_1_15_port, A1 => n143, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_15_port, 
                           B1 => input_previous_1_17_port, Y => n4434);
   U6181 : XNOR2X1 port map( A => n3689, B => input_previous_1_15_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_15_port);
   U6182 : AOI22X1 port map( A0 => input_previous_0_15_port, A1 => n131, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_15_port, 
                           B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn83);
   U6183 : XNOR2X1 port map( A => n3641, B => input_previous_0_15_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_15_port);
   U6184 : INVX1 port map( A => input_previous_1_17_port, Y => n254);
   U6185 : INVX1 port map( A => input_previous_2_17_port, Y => n255);
   U6186 : INVX1 port map( A => output_previous_2_17_port, Y => n256);
   U6187 : INVX1 port map( A => input_previous_0_17_port, Y => n282);
   U6188 : BUFX3 port map( A => n4478, Y => n202);
   U6189 : AOI22X1 port map( A0 => input_previous_2_8_port, A1 => n142, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_8_port, 
                           B1 => input_previous_2_17_port, Y => n4478);
   U6190 : XOR2X1 port map( A => n3728, B => input_previous_2_8_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_8_port);
   U6191 : OR2X2 port map( A => input_previous_2_7_port, B => n3729, Y => n3728
                           );
   U6192 : BUFX3 port map( A => n4584, Y => n244);
   U6193 : AOI22X1 port map( A0 => output_previous_2_8_port, A1 => n140, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_8_port, 
                           B1 => output_previous_2_17_port, Y => n4584);
   U6194 : XOR2X1 port map( A => n3824, B => output_previous_2_8_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_8_port);
   U6195 : OR2X2 port map( A => output_previous_2_7_port, B => n3825, Y => 
                           n3824);
   U6196 : BUFX3 port map( A => n4483, Y => n207);
   U6197 : AOI22X1 port map( A0 => input_previous_2_3_port, A1 => n142, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_3_port, 
                           B1 => input_previous_2_17_port, Y => n4483);
   U6198 : XOR2X1 port map( A => n3733, B => input_previous_2_3_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_3_port);
   U6199 : BUFX3 port map( A => n4589, Y => n249);
   U6200 : AOI22X1 port map( A0 => output_previous_2_3_port, A1 => n140, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_3_port, 
                           B1 => output_previous_2_17_port, Y => n4589);
   U6201 : XOR2X1 port map( A => n3829, B => output_previous_2_3_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_3_port);
   U6202 : AOI22X1 port map( A0 => input_previous_1_12_port, A1 => n143, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_12_port, 
                           B1 => input_previous_1_17_port, Y => n4437);
   U6203 : XOR2X1 port map( A => n3693, B => input_previous_1_12_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_12_port);
   U6204 : OR2X2 port map( A => n3692, B => input_previous_1_11_port, Y => 
                           n3693);
   U6205 : AOI22X1 port map( A0 => input_previous_0_12_port, A1 => n131, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_12_port, 
                           B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn86);
   U6206 : XOR2X1 port map( A => n3645, B => input_previous_0_12_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_12_port);
   U6207 : OR2X2 port map( A => n3644, B => input_previous_0_11_port, Y => 
                           n3645);
   U6208 : BUFX3 port map( A => n4425, Y => n181);
   U6209 : AOI22X1 port map( A0 => input_previous_1_8_port, A1 => n144, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_8_port, 
                           B1 => input_previous_1_17_port, Y => n4425);
   U6210 : XOR2X1 port map( A => n3680, B => input_previous_1_8_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_8_port);
   U6211 : OR2X2 port map( A => input_previous_1_7_port, B => n3681, Y => n3680
                           );
   U6212 : BUFX3 port map( A => input_times_b0_mul_componentxn74, Y => n272);
   U6213 : AOI22X1 port map( A0 => input_previous_0_8_port, A1 => n132, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_8_port
                           , B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn74);
   U6214 : XOR2X1 port map( A => n3632, B => input_previous_0_8_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_8_port
                           );
   U6215 : OR2X2 port map( A => input_previous_0_7_port, B => n3633, Y => n3632
                           );
   U6216 : BUFX3 port map( A => n4482, Y => n206);
   U6217 : AOI22X1 port map( A0 => input_previous_2_4_port, A1 => n142, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_4_port, 
                           B1 => input_previous_2_17_port, Y => n4482);
   U6218 : XOR2X1 port map( A => n3732, B => input_previous_2_4_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_4_port);
   U6219 : OR2X2 port map( A => input_previous_2_3_port, B => n3733, Y => n3732
                           );
   U6220 : BUFX3 port map( A => n4588, Y => n248);
   U6221 : AOI22X1 port map( A0 => output_previous_2_4_port, A1 => n140, B0 => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_4_port, 
                           B1 => output_previous_2_17_port, Y => n4588);
   U6222 : XOR2X1 port map( A => n3828, B => output_previous_2_4_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_4_port);
   U6223 : OR2X2 port map( A => output_previous_2_3_port, B => n3829, Y => 
                           n3828);
   U6224 : AOI22X1 port map( A0 => input_previous_1_16_port, A1 => n143, B0 => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_16_port, 
                           B1 => input_previous_1_17_port, Y => n4433);
   U6225 : XNOR2X1 port map( A => n3688, B => input_previous_1_16_port, Y => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_16_port);
   U6226 : AOI22X1 port map( A0 => input_previous_2_16_port, A1 => n141, B0 => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_16_port, 
                           B1 => input_previous_2_17_port, Y => n4486);
   U6227 : XNOR2X1 port map( A => n3736, B => input_previous_2_16_port, Y => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_16_port);
   U6228 : AOI22X1 port map( A0 => output_previous_2_16_port, A1 => n139, B0 =>
                           output_p2_times_a2_mul_componentxinput_A_inverted_16_port, 
                           B1 => output_previous_2_17_port, Y => n4592);
   U6229 : XNOR2X1 port map( A => n3832, B => output_previous_2_16_port, Y => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_16_port);
   U6230 : AOI22X1 port map( A0 => input_previous_0_16_port, A1 => n131, B0 => 
                           input_times_b0_mul_componentxinput_A_inverted_16_port, 
                           B1 => input_previous_0_17_port, Y => 
                           input_times_b0_mul_componentxn82);
   U6231 : XNOR2X1 port map( A => n3640, B => input_previous_0_16_port, Y => 
                           input_times_b0_mul_componentxinput_A_inverted_16_port);
   U6232 : NOR2BX1 port map( AN => n3689, B => input_previous_1_15_port, Y => 
                           n3688);
   U6233 : NOR2BX1 port map( AN => n3641, B => input_previous_0_15_port, Y => 
                           n3640);
   U6234 : NOR2BX1 port map( AN => n3737, B => input_previous_2_15_port, Y => 
                           n3736);
   U6235 : NOR2BX1 port map( AN => n3833, B => output_previous_2_15_port, Y => 
                           n3832);
   U6236 : INVX1 port map( A => input_previous_1_9_port, Y => n1293);
   U6237 : INVX1 port map( A => input_previous_0_9_port, Y => n1191);
   U6238 : NAND2BX1 port map( AN => input_previous_1_16_port, B => n3688, Y => 
                           n3687);
   U6239 : NAND2BX1 port map( AN => input_previous_0_16_port, B => n3640, Y => 
                           n3639);
   U6240 : NAND2BX1 port map( AN => input_previous_2_16_port, B => n3736, Y => 
                           n3735);
   U6241 : NAND2BX1 port map( AN => output_previous_2_16_port, B => n3832, Y =>
                           n3831);
   U6242 : INVX1 port map( A => input_previous_2_9_port, Y => n1283);
   U6243 : INVX1 port map( A => output_previous_2_9_port, Y => n1282);
   U6244 : OAI2BB2X1 port map( B0 => n1214, B1 => n1260, A0N => 
                           output_previous_2_7_port, A1N => n320, Y => n4662);
   U6245 : INVX1 port map( A => output_signal_7_port, Y => n1214);
   U6246 : OAI2BB2X1 port map( B0 => n1218, B1 => n321, A0N => 
                           output_previous_2_5_port, A1N => n320, Y => n4660);
   U6247 : INVX1 port map( A => output_signal_5_port, Y => n1218);
   U6248 : OAI2BB2X1 port map( B0 => n1216, B1 => n1260, A0N => 
                           output_previous_2_6_port, A1N => n320, Y => n4661);
   U6249 : INVX1 port map( A => output_signal_6_port, Y => n1216);
   U6250 : OAI2BB2X1 port map( B0 => n1202, B1 => n1260, A0N => 
                           output_previous_2_15_port, A1N => n319, Y => n4670);
   U6251 : INVX1 port map( A => output_previous_1_15_port, Y => n1202);
   U6252 : OAI2BB2X1 port map( B0 => n1201, B1 => n320, A0N => 
                           output_previous_2_14_port, A1N => n319, Y => n4669);
   U6253 : INVX1 port map( A => output_previous_1_14_port, Y => n1201);
   U6254 : OAI2BB2X1 port map( B0 => n1200, B1 => n319, A0N => 
                           output_previous_2_13_port, A1N => n319, Y => n4668);
   U6255 : INVX1 port map( A => output_previous_1_13_port, Y => n1200);
   U6256 : OAI2BB2X1 port map( B0 => n1204, B1 => n1260, A0N => 
                           output_previous_2_16_port, A1N => n319, Y => n4671);
   U6257 : INVX1 port map( A => output_previous_1_16_port, Y => n1204);
   U6258 : OAI2BB2X1 port map( B0 => n1224, B1 => n1260, A0N => 
                           output_previous_2_2_port, A1N => n320, Y => n4657);
   U6259 : INVX1 port map( A => output_signal_2_port, Y => n1224);
   U6260 : OAI2BB2X1 port map( B0 => n1222, B1 => n319, A0N => 
                           output_previous_2_3_port, A1N => n320, Y => n4658);
   U6261 : INVX1 port map( A => output_signal_3_port, Y => n1222);
   U6262 : OAI2BB2X1 port map( B0 => n1220, B1 => n1260, A0N => 
                           output_previous_2_4_port, A1N => n320, Y => n4659);
   U6263 : INVX1 port map( A => output_signal_4_port, Y => n1220);
   U6264 : OAI2BB2X1 port map( B0 => n1206, B1 => n319, A0N => 
                           output_previous_2_11_port, A1N => n320, Y => n4666);
   U6265 : INVX1 port map( A => output_previous_1_11_port, Y => n1206);
   U6266 : OAI2BB2X1 port map( B0 => n1208, B1 => n1260, A0N => 
                           output_previous_2_10_port, A1N => n320, Y => n4665);
   U6267 : INVX1 port map( A => output_previous_1_10_port, Y => n1208);
   U6268 : OAI2BB2X1 port map( B0 => n1210, B1 => n321, A0N => 
                           output_previous_2_9_port, A1N => n320, Y => n4664);
   U6269 : OAI2BB2X1 port map( B0 => n1199, B1 => n1260, A0N => 
                           output_previous_2_12_port, A1N => n320, Y => n4667);
   U6270 : INVX1 port map( A => output_previous_1_12_port, Y => n1199);
   U6271 : AOI32X1 port map( A0 => n846, A1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn18, 
                           A2 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_0, 
                           B0 => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_1_port, 
                           B1 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_1, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn16);
   U6272 : AOI32X1 port map( A0 => n1005, A1 => n1650, A2 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_0, 
                           B0 => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_1_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1648);
   U6273 : AOI32X1 port map( A0 => n1164, A1 => n1682, A2 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_0, 
                           B0 => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_1_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1680);
   U6274 : AOI32X1 port map( A0 => n528, A1 => n1714, A2 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_0, 
                           B0 => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_1_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1712);
   U6275 : AOI32X1 port map( A0 => n687, A1 => n1746, A2 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_0, 
                           B0 => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_1_port, 
                           B1 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1744);
   U6276 : OAI221XL port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_8, 
                           A1 => input_times_b0_div_componentxn53, B0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_9, 
                           B1 => input_times_b0_div_componentxn54, C0 => n1546,
                           Y => n1547);
   U6277 : OAI221XL port map( A0 => n853, A1 => n1531, B0 => n854, B1 => n1530,
                           C0 => n1545, Y => n1546);
   U6278 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1530);
   U6279 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_7, Y 
                           => n1531);
   U6280 : OAI221XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n4231, B0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_9, 
                           B1 => n4232, C0 => n1622, Y => n1623);
   U6281 : OAI221XL port map( A0 => n1012, A1 => n1515, B0 => n1013, B1 => 
                           n1514, C0 => n1621, Y => n1622);
   U6282 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1514);
   U6283 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_7, Y 
                           => n1515);
   U6284 : OAI221XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n4287, B0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_9, 
                           B1 => n4288, C0 => n1603, Y => n1604);
   U6285 : OAI221XL port map( A0 => n1171, A1 => n1499, B0 => n1172, B1 => 
                           n1498, C0 => n1602, Y => n1603);
   U6286 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1498);
   U6287 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_7, Y 
                           => n1499);
   U6288 : OAI221XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n4341, B0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_9, 
                           B1 => n4342, C0 => n1584, Y => n1585);
   U6289 : OAI221XL port map( A0 => n535, A1 => n1483, B0 => n536, B1 => n1482,
                           C0 => n1583, Y => n1584);
   U6290 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1482);
   U6291 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_7, Y 
                           => n1483);
   U6292 : OAI221XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n4397, B0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_9, 
                           B1 => n4398, C0 => n1565, Y => n1566);
   U6293 : OAI221XL port map( A0 => n694, A1 => n1467, B0 => n695, B1 => n1466,
                           C0 => n1564, Y => n1565);
   U6294 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1466);
   U6295 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_7, Y 
                           => n1467);
   U6296 : OAI221XL port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_2, 
                           A1 => input_times_b0_div_componentxn47, B0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_3, 
                           B1 => input_times_b0_div_componentxn48, C0 => n1540,
                           Y => n1541);
   U6297 : OAI222XL port map( A0 => n1539, A1 => n1537, B0 => n847, B1 => n1538
                           , C0 => n848, C1 => n1536, Y => n1540);
   U6298 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1536);
   U6299 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1537);
   U6300 : OAI221XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n4225, B0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_3, 
                           B1 => n4226, C0 => n1616, Y => n1617);
   U6301 : OAI222XL port map( A0 => n1615, A1 => n1521, B0 => n1006, B1 => 
                           n1614, C0 => n1007, C1 => n1520, Y => n1616);
   U6302 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1520);
   U6303 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1521);
   U6304 : OAI221XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n4281, B0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_3, 
                           B1 => n4282, C0 => n1597, Y => n1598);
   U6305 : OAI222XL port map( A0 => n1596, A1 => n1505, B0 => n1165, B1 => 
                           n1595, C0 => n1166, C1 => n1504, Y => n1597);
   U6306 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1504);
   U6307 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1505);
   U6308 : OAI221XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n4335, B0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_3, 
                           B1 => n4336, C0 => n1578, Y => n1579);
   U6309 : OAI222XL port map( A0 => n1577, A1 => n1489, B0 => n529, B1 => n1576
                           , C0 => n530, C1 => n1488, Y => n1578);
   U6310 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1488);
   U6311 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1489);
   U6312 : OAI221XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n4391, B0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_3, 
                           B1 => n4392, C0 => n1559, Y => n1560);
   U6313 : OAI222XL port map( A0 => n1558, A1 => n1473, B0 => n688, B1 => n1557
                           , C0 => n689, C1 => n1472, Y => n1559);
   U6314 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1472);
   U6315 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1473);
   U6316 : OAI221XL port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_4, 
                           A1 => input_times_b0_div_componentxn49, B0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_5, 
                           B1 => input_times_b0_div_componentxn50, C0 => n1542,
                           Y => n1543);
   U6317 : OAI221XL port map( A0 => n849, A1 => n1535, B0 => n850, B1 => n1534,
                           C0 => n1541, Y => n1542);
   U6318 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1534);
   U6319 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_3, Y 
                           => n1535);
   U6320 : OAI221XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n4227, B0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_5, 
                           B1 => n4228, C0 => n1618, Y => n1619);
   U6321 : OAI221XL port map( A0 => n1008, A1 => n1519, B0 => n1009, B1 => 
                           n1518, C0 => n1617, Y => n1618);
   U6322 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1518);
   U6323 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_3, Y 
                           => n1519);
   U6324 : OAI221XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n4283, B0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_5, 
                           B1 => n4284, C0 => n1599, Y => n1600);
   U6325 : OAI221XL port map( A0 => n1167, A1 => n1503, B0 => n1168, B1 => 
                           n1502, C0 => n1598, Y => n1599);
   U6326 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1502);
   U6327 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_3, Y 
                           => n1503);
   U6328 : OAI221XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n4337, B0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_5, 
                           B1 => n4338, C0 => n1580, Y => n1581);
   U6329 : OAI221XL port map( A0 => n531, A1 => n1487, B0 => n532, B1 => n1486,
                           C0 => n1579, Y => n1580);
   U6330 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1486);
   U6331 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_3, Y 
                           => n1487);
   U6332 : OAI221XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n4393, B0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_5, 
                           B1 => n4394, C0 => n1561, Y => n1562);
   U6333 : OAI221XL port map( A0 => n690, A1 => n1471, B0 => n691, B1 => n1470,
                           C0 => n1560, Y => n1561);
   U6334 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1470);
   U6335 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_3, Y 
                           => n1471);
   U6336 : OAI221XL port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_6, 
                           A1 => input_times_b0_div_componentxn51, B0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_7, 
                           B1 => input_times_b0_div_componentxn52, C0 => n1544,
                           Y => n1545);
   U6337 : OAI221XL port map( A0 => n851, A1 => n1533, B0 => n852, B1 => n1532,
                           C0 => n1543, Y => n1544);
   U6338 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1532);
   U6339 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_5, Y 
                           => n1533);
   U6340 : OAI221XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n4229, B0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_7, 
                           B1 => n4230, C0 => n1620, Y => n1621);
   U6341 : OAI221XL port map( A0 => n1010, A1 => n1517, B0 => n1011, B1 => 
                           n1516, C0 => n1619, Y => n1620);
   U6342 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1516);
   U6343 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_5, Y 
                           => n1517);
   U6344 : OAI221XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n4285, B0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_7, 
                           B1 => n4286, C0 => n1601, Y => n1602);
   U6345 : OAI221XL port map( A0 => n1169, A1 => n1501, B0 => n1170, B1 => 
                           n1500, C0 => n1600, Y => n1601);
   U6346 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1500);
   U6347 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_5, Y 
                           => n1501);
   U6348 : OAI221XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n4339, B0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_7, 
                           B1 => n4340, C0 => n1582, Y => n1583);
   U6349 : OAI221XL port map( A0 => n533, A1 => n1485, B0 => n534, B1 => n1484,
                           C0 => n1581, Y => n1582);
   U6350 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1484);
   U6351 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_5, Y 
                           => n1485);
   U6352 : OAI221XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n4395, B0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_7, 
                           B1 => n4396, C0 => n1563, Y => n1564);
   U6353 : OAI221XL port map( A0 => n692, A1 => n1469, B0 => n693, B1 => n1468,
                           C0 => n1562, Y => n1563);
   U6354 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1468);
   U6355 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_5, Y 
                           => n1469);
   U6356 : OAI221XL port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_10, 
                           A1 => input_times_b0_div_componentxn55, B0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_11, 
                           B1 => input_times_b0_div_componentxn56, C0 => n1548,
                           Y => n1549);
   U6357 : OAI221XL port map( A0 => n845, A1 => n1528, B0 => n855, B1 => n1529,
                           C0 => n1547, Y => n1548);
   U6358 : INVX1 port map( A => input_times_b0_div_componentxn54, Y => n855);
   U6359 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1528);
   U6360 : OAI221XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n4233, B0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_11, 
                           B1 => n4234, C0 => n1624, Y => n1625);
   U6361 : OAI221XL port map( A0 => n1004, A1 => n1512, B0 => n1014, B1 => 
                           n1513, C0 => n1623, Y => n1624);
   U6362 : INVX1 port map( A => n4232, Y => n1014);
   U6363 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1512);
   U6364 : OAI221XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n4289, B0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_11, 
                           B1 => n4290, C0 => n1605, Y => n1606);
   U6365 : OAI221XL port map( A0 => n1163, A1 => n1496, B0 => n1173, B1 => 
                           n1497, C0 => n1604, Y => n1605);
   U6366 : INVX1 port map( A => n4288, Y => n1173);
   U6367 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1496);
   U6368 : OAI221XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n4343, B0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_11, 
                           B1 => n4344, C0 => n1586, Y => n1587);
   U6369 : OAI221XL port map( A0 => n527, A1 => n1480, B0 => n537, B1 => n1481,
                           C0 => n1585, Y => n1586);
   U6370 : INVX1 port map( A => n4342, Y => n537);
   U6371 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1480);
   U6372 : OAI221XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n4399, B0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_11, 
                           B1 => n4400, C0 => n1567, Y => n1568);
   U6373 : OAI221XL port map( A0 => n686, A1 => n1464, B0 => n696, B1 => n1465,
                           C0 => n1566, Y => n1567);
   U6374 : INVX1 port map( A => n4398, Y => n696);
   U6375 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1464);
   U6376 : OAI221XL port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_12, 
                           A1 => input_times_b0_div_componentxn57, B0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_13, 
                           B1 => input_times_b0_div_componentxn58, C0 => n1550,
                           Y => n1551);
   U6377 : OAI221XL port map( A0 => n838, A1 => n1527, B0 => n839, B1 => n1526,
                           C0 => n1549, Y => n1550);
   U6378 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1526);
   U6379 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_11, Y 
                           => n1527);
   U6380 : OAI221XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n4235, B0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_13, 
                           B1 => n4236, C0 => n1626, Y => n1627);
   U6381 : OAI221XL port map( A0 => n997, A1 => n1511, B0 => n998, B1 => n1510,
                           C0 => n1625, Y => n1626);
   U6382 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1510);
   U6383 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_11, Y 
                           => n1511);
   U6384 : OAI221XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n4291, B0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_13, 
                           B1 => n4292, C0 => n1607, Y => n1608);
   U6385 : OAI221XL port map( A0 => n1156, A1 => n1495, B0 => n1157, B1 => 
                           n1494, C0 => n1606, Y => n1607);
   U6386 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1494);
   U6387 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_11, Y 
                           => n1495);
   U6388 : OAI221XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n4345, B0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_13, 
                           B1 => n4346, C0 => n1588, Y => n1589);
   U6389 : OAI221XL port map( A0 => n520, A1 => n1479, B0 => n521, B1 => n1478,
                           C0 => n1587, Y => n1588);
   U6390 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1478);
   U6391 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_11, Y 
                           => n1479);
   U6392 : OAI221XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n4401, B0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_13, 
                           B1 => n4402, C0 => n1569, Y => n1570);
   U6393 : OAI221XL port map( A0 => n679, A1 => n1463, B0 => n680, B1 => n1462,
                           C0 => n1568, Y => n1569);
   U6394 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1462);
   U6395 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_11, Y 
                           => n1463);
   U6396 : OAI221XL port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_14, 
                           A1 => input_times_b0_div_componentxn59, B0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_15, 
                           B1 => input_times_b0_div_componentxn60, C0 => n1552,
                           Y => n1553);
   U6397 : OAI221XL port map( A0 => n840, A1 => n1525, B0 => n841, B1 => n1524,
                           C0 => n1551, Y => n1552);
   U6398 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1524);
   U6399 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_13, Y 
                           => n1525);
   U6400 : OAI221XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n4237, B0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_15, 
                           B1 => n4238, C0 => n1628, Y => n1629);
   U6401 : OAI221XL port map( A0 => n999, A1 => n1509, B0 => n1000, B1 => n1508
                           , C0 => n1627, Y => n1628);
   U6402 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1508);
   U6403 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_13, Y 
                           => n1509);
   U6404 : OAI221XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n4293, B0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_15, 
                           B1 => n4294, C0 => n1609, Y => n1610);
   U6405 : OAI221XL port map( A0 => n1158, A1 => n1493, B0 => n1159, B1 => 
                           n1492, C0 => n1608, Y => n1609);
   U6406 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1492);
   U6407 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_13, Y 
                           => n1493);
   U6408 : OAI221XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n4347, B0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_15, 
                           B1 => n4348, C0 => n1590, Y => n1591);
   U6409 : OAI221XL port map( A0 => n522, A1 => n1477, B0 => n523, B1 => n1476,
                           C0 => n1589, Y => n1590);
   U6410 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1476);
   U6411 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_13, Y 
                           => n1477);
   U6412 : OAI221XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n4403, B0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_15, 
                           B1 => n4404, C0 => n1571, Y => n1572);
   U6413 : OAI221XL port map( A0 => n681, A1 => n1461, B0 => n682, B1 => n1460,
                           C0 => n1570, Y => n1571);
   U6414 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1460);
   U6415 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_13, Y 
                           => n1461);
   U6416 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_3_port, 
                           A1 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_3, 
                           B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn13, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn14, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn12);
   U6417 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_3_port, 
                           A1 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n1645, B1 => n1646, Y => n1644);
   U6418 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_3_port, 
                           A1 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n1677, B1 => n1678, Y => n1676);
   U6419 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_3_port, 
                           A1 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n1709, B1 => n1710, Y => n1708);
   U6420 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_3_port, 
                           A1 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n1741, B1 => n1742, Y => n1740);
   U6421 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_5_port, 
                           A1 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_5, 
                           B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn9, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn10, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn8);
   U6422 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_5_port, 
                           A1 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n1641, B1 => n1642, Y => n1640);
   U6423 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_5_port, 
                           A1 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n1673, B1 => n1674, Y => n1672);
   U6424 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_5_port, 
                           A1 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n1705, B1 => n1706, Y => n1704);
   U6425 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_5_port, 
                           A1 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n1737, B1 => n1738, Y => n1736);
   U6426 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_7_port, 
                           A1 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_7, 
                           B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn5, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn6, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn4);
   U6427 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_7_port, 
                           A1 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n1637, B1 => n1638, Y => n1636);
   U6428 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_7_port, 
                           A1 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n1669, B1 => n1670, Y => n1668);
   U6429 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_7_port, 
                           A1 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n1701, B1 => n1702, Y => n1700);
   U6430 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_7_port, 
                           A1 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n1733, B1 => n1734, Y => n1732);
   U6431 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_9_port, 
                           A1 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_9, 
                           B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn1, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn2, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn35);
   U6432 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_9_port, 
                           A1 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n1633, B1 => n1634, Y => n1663);
   U6433 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_9_port, 
                           A1 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n1665, B1 => n1666, Y => n1695);
   U6434 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_9_port, 
                           A1 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n1697, B1 => n1698, Y => n1727);
   U6435 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_9_port, 
                           A1 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n1729, B1 => n1730, Y => n1759);
   U6436 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_11_port, 
                           A1 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_11, 
                           B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn33, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn34, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn31);
   U6437 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_11_port, 
                           A1 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n1661, B1 => n1662, Y => n1659);
   U6438 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_11_port, 
                           A1 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n1693, B1 => n1694, Y => n1691);
   U6439 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_11_port, 
                           A1 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n1725, B1 => n1726, Y => n1723);
   U6440 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_11_port, 
                           A1 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n1757, B1 => n1758, Y => n1755);
   U6441 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_13_port, 
                           A1 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_13, 
                           B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn29, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn30, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn27);
   U6442 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_13_port, 
                           A1 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n1657, B1 => n1658, Y => n1655);
   U6443 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_13_port, 
                           A1 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n1689, B1 => n1690, Y => n1687);
   U6444 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_13_port, 
                           A1 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n1721, B1 => n1722, Y => n1719);
   U6445 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_13_port, 
                           A1 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n1753, B1 => n1754, Y => n1751);
   U6446 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn16, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn15, 
                           A0N => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_2_port, 
                           A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_2, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn13);
   U6447 : OAI2BB2X1 port map( B0 => n1648, B1 => n1647, A0N => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_2_port, 
                           A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1645);
   U6448 : OAI2BB2X1 port map( B0 => n1680, B1 => n1679, A0N => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_2_port, 
                           A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1677);
   U6449 : OAI2BB2X1 port map( B0 => n1712, B1 => n1711, A0N => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_2_port, 
                           A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1709);
   U6450 : OAI2BB2X1 port map( B0 => n1744, B1 => n1743, A0N => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_2_port, 
                           A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_2, Y 
                           => n1741);
   U6451 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn12, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn11, 
                           A0N => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_4_port, 
                           A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_4, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn9);
   U6452 : OAI2BB2X1 port map( B0 => n1644, B1 => n1643, A0N => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_4_port, 
                           A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1641);
   U6453 : OAI2BB2X1 port map( B0 => n1676, B1 => n1675, A0N => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_4_port, 
                           A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1673);
   U6454 : OAI2BB2X1 port map( B0 => n1708, B1 => n1707, A0N => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_4_port, 
                           A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1705);
   U6455 : OAI2BB2X1 port map( B0 => n1740, B1 => n1739, A0N => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_4_port, 
                           A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_4, Y 
                           => n1737);
   U6456 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn8, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn7, 
                           A0N => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_6_port, 
                           A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_6, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn5);
   U6457 : OAI2BB2X1 port map( B0 => n1640, B1 => n1639, A0N => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_6_port, 
                           A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1637);
   U6458 : OAI2BB2X1 port map( B0 => n1672, B1 => n1671, A0N => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_6_port, 
                           A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1669);
   U6459 : OAI2BB2X1 port map( B0 => n1704, B1 => n1703, A0N => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_6_port, 
                           A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1701);
   U6460 : OAI2BB2X1 port map( B0 => n1736, B1 => n1735, A0N => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_6_port, 
                           A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_6, Y 
                           => n1733);
   U6461 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn4, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn3, 
                           A0N => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_8_port, 
                           A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_8, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn1);
   U6462 : OAI2BB2X1 port map( B0 => n1636, B1 => n1635, A0N => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_8_port, 
                           A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1633);
   U6463 : OAI2BB2X1 port map( B0 => n1668, B1 => n1667, A0N => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_8_port, 
                           A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1665);
   U6464 : OAI2BB2X1 port map( B0 => n1700, B1 => n1699, A0N => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_8_port, 
                           A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1697);
   U6465 : OAI2BB2X1 port map( B0 => n1732, B1 => n1731, A0N => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_8_port, 
                           A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_8, Y 
                           => n1729);
   U6466 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn35, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn36, 
                           A0N => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_10_port, 
                           A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_10, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn33);
   U6467 : OAI2BB2X1 port map( B0 => n1663, B1 => n1664, A0N => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_10_port, 
                           A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1661);
   U6468 : OAI2BB2X1 port map( B0 => n1695, B1 => n1696, A0N => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_10_port, 
                           A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1693);
   U6469 : OAI2BB2X1 port map( B0 => n1727, B1 => n1728, A0N => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_10_port, 
                           A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1725);
   U6470 : OAI2BB2X1 port map( B0 => n1759, B1 => n1760, A0N => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_10_port, 
                           A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_10, Y 
                           => n1757);
   U6471 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn31, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn32, 
                           A0N => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_12_port, 
                           A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_12, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn29);
   U6472 : OAI2BB2X1 port map( B0 => n1659, B1 => n1660, A0N => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_12_port, 
                           A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1657);
   U6473 : OAI2BB2X1 port map( B0 => n1691, B1 => n1692, A0N => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_12_port, 
                           A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1689);
   U6474 : OAI2BB2X1 port map( B0 => n1723, B1 => n1724, A0N => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_12_port, 
                           A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1721);
   U6475 : OAI2BB2X1 port map( B0 => n1755, B1 => n1756, A0N => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_12_port, 
                           A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_12, Y 
                           => n1753);
   U6476 : OAI2BB2X1 port map( B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn27, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn28, 
                           A0N => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_14_port, 
                           A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_14, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn25);
   U6477 : OAI2BB2X1 port map( B0 => n1655, B1 => n1656, A0N => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_14_port, 
                           A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1653);
   U6478 : OAI2BB2X1 port map( B0 => n1687, B1 => n1688, A0N => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_14_port, 
                           A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1685);
   U6479 : OAI2BB2X1 port map( B0 => n1719, B1 => n1720, A0N => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_14_port, 
                           A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1717);
   U6480 : OAI2BB2X1 port map( B0 => n1751, B1 => n1752, A0N => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_14_port, 
                           A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_14, Y 
                           => n1749);
   U6481 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_15_port, 
                           A1 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_15, 
                           B0 => 
                           input_times_b0_div_componentxUDxactually_substractsxn25, 
                           B1 => 
                           input_times_b0_div_componentxUDxactually_substractsxn26, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn23);
   U6482 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_15_port, 
                           A1 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n1653, B1 => n1654, Y => n1651);
   U6483 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_15_port, 
                           A1 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n1685, B1 => n1686, Y => n1683);
   U6484 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_15_port, 
                           A1 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n1717, B1 => n1718, Y => n1715);
   U6485 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_15_port, 
                           A1 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n1749, B1 => n1750, Y => n1747);
   U6486 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_3, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_3_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn14);
   U6487 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_3, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_3_port, Y 
                           => n1646);
   U6488 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_3, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_3_port, Y 
                           => n1678);
   U6489 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_3, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_3_port, Y 
                           => n1710);
   U6490 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_3, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_3_port, Y 
                           => n1742);
   U6491 : NOR2BX1 port map( AN => n846, B => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_0, Y 
                           => n1539);
   U6492 : NOR2BX1 port map( AN => n1005, B => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_0, Y 
                           => n1615);
   U6493 : NOR2BX1 port map( AN => n1164, B => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_0, Y 
                           => n1596);
   U6494 : NOR2BX1 port map( AN => n528, B => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_0, Y 
                           => n1577);
   U6495 : NOR2BX1 port map( AN => n687, B => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_0, Y 
                           => n1558);
   U6496 : OAI2BB2X1 port map( B0 => n1236, B1 => n1260, A0N => 
                           output_p2_times_a2_mul_componentxinput_A_inverted_0_port, 
                           A1N => n320, Y => n4655);
   U6497 : INVX1 port map( A => 
                           output_p1_times_a1_mul_componentxinput_A_inverted_0_port, Y 
                           => n1236);
   U6498 : OAI2BB2X1 port map( B0 => n1226, B1 => n1260, A0N => 
                           output_previous_2_1_port, A1N => n320, Y => n4656);
   U6499 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_1, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_1_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn18);
   U6500 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_1, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_1_port, Y 
                           => n1650);
   U6501 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_1, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_1_port, Y 
                           => n1682);
   U6502 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_1, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_1_port, Y 
                           => n1714);
   U6503 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_1, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_1_port, Y 
                           => n1746);
   U6504 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_2, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_2_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn15);
   U6505 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_2, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_2_port, Y 
                           => n1647);
   U6506 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_2, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_2_port, Y 
                           => n1679);
   U6507 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_2, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_2_port, Y 
                           => n1711);
   U6508 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_2, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_2_port, Y 
                           => n1743);
   U6509 : OAI2BB2X1 port map( B0 => n1212, B1 => n320, A0N => 
                           output_previous_2_8_port, A1N => n320, Y => n4663);
   U6510 : INVX1 port map( A => output_previous_1_8_port, Y => n1212);
   U6511 : NOR2BX1 port map( AN => n1539, B => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1538);
   U6512 : NOR2BX1 port map( AN => n1615, B => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1614);
   U6513 : NOR2BX1 port map( AN => n1596, B => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1595);
   U6514 : NOR2BX1 port map( AN => n1577, B => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1576);
   U6515 : NOR2BX1 port map( AN => n1558, B => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_1, Y 
                           => n1557);
   U6516 : OAI2BB1X1 port map( A0N => n1522, A1N => n843, B0 => n1554, Y => 
                           n1555);
   U6517 : OAI221XL port map( A0 => n842, A1 => n1523, B0 => n843, B1 => n1522,
                           C0 => n1553, Y => n1554);
   U6518 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_16, Y 
                           => n1522);
   U6519 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_15, Y 
                           => n1523);
   U6520 : OAI2BB1X1 port map( A0N => n1506, A1N => n1002, B0 => n1630, Y => 
                           n1631);
   U6521 : OAI221XL port map( A0 => n1001, A1 => n1507, B0 => n1002, B1 => 
                           n1506, C0 => n1629, Y => n1630);
   U6522 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_16, Y 
                           => n1506);
   U6523 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_15, Y 
                           => n1507);
   U6524 : OAI2BB1X1 port map( A0N => n1490, A1N => n1161, B0 => n1611, Y => 
                           n1612);
   U6525 : OAI221XL port map( A0 => n1160, A1 => n1491, B0 => n1161, B1 => 
                           n1490, C0 => n1610, Y => n1611);
   U6526 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_16, Y 
                           => n1490);
   U6527 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_15, Y 
                           => n1491);
   U6528 : OAI2BB1X1 port map( A0N => n1474, A1N => n525, B0 => n1592, Y => 
                           n1593);
   U6529 : OAI221XL port map( A0 => n524, A1 => n1475, B0 => n525, B1 => n1474,
                           C0 => n1591, Y => n1592);
   U6530 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_16, Y 
                           => n1474);
   U6531 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_15, Y 
                           => n1475);
   U6532 : OAI2BB1X1 port map( A0N => n1458, A1N => n684, B0 => n1573, Y => 
                           n1574);
   U6533 : OAI221XL port map( A0 => n683, A1 => n1459, B0 => n684, B1 => n1458,
                           C0 => n1572, Y => n1573);
   U6534 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_16, Y 
                           => n1458);
   U6535 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_15, Y 
                           => n1459);
   U6536 : INVX1 port map( A => input_times_b0_div_componentxUDxis_less_than, Y
                           => n837);
   U6537 : OAI21XL port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_17, 
                           A1 => n844, B0 => n1556, Y => 
                           input_times_b0_div_componentxUDxis_less_than);
   U6538 : OAI2BB1X1 port map( A0N => n844, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_17, 
                           B0 => n1555, Y => n1556);
   U6539 : INVX1 port map( A => input_times_b0_div_componentxunsigned_B_17, Y 
                           => n844);
   U6540 : INVX1 port map( A => input_p1_times_b1_div_componentxUDxis_less_than
                           , Y => n996);
   U6541 : OAI21XL port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_17, 
                           A1 => n1003, B0 => n1632, Y => 
                           input_p1_times_b1_div_componentxUDxis_less_than);
   U6542 : OAI2BB1X1 port map( A0N => n1003, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_17, 
                           B0 => n1631, Y => n1632);
   U6543 : INVX1 port map( A => input_p1_times_b1_div_componentxunsigned_B_17, 
                           Y => n1003);
   U6544 : INVX1 port map( A => input_p2_times_b2_div_componentxUDxis_less_than
                           , Y => n1155);
   U6545 : OAI21XL port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_17, 
                           A1 => n1162, B0 => n1613, Y => 
                           input_p2_times_b2_div_componentxUDxis_less_than);
   U6546 : OAI2BB1X1 port map( A0N => n1162, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_17, 
                           B0 => n1612, Y => n1613);
   U6547 : INVX1 port map( A => input_p2_times_b2_div_componentxunsigned_B_17, 
                           Y => n1162);
   U6548 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxis_less_than, Y 
                           => n519);
   U6549 : OAI21XL port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_17, 
                           A1 => n526, B0 => n1594, Y => 
                           output_p1_times_a1_div_componentxUDxis_less_than);
   U6550 : OAI2BB1X1 port map( A0N => n526, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_17, 
                           B0 => n1593, Y => n1594);
   U6551 : INVX1 port map( A => output_p1_times_a1_div_componentxunsigned_B_17,
                           Y => n526);
   U6552 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxis_less_than, Y 
                           => n678);
   U6553 : OAI21XL port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_17, 
                           A1 => n685, B0 => n1575, Y => 
                           output_p2_times_a2_div_componentxUDxis_less_than);
   U6554 : OAI2BB1X1 port map( A0N => n685, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_17, 
                           B0 => n1574, Y => n1575);
   U6555 : INVX1 port map( A => output_p2_times_a2_div_componentxunsigned_B_17,
                           Y => n685);
   U6556 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_4, 
                           B0 => n1810, Y => n1828);
   U6557 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_3, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_3_port, 
                           B1 => n14, Y => n1810);
   U6558 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn13, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn14, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_3_port);
   U6559 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_6, 
                           B0 => n1808, Y => n1826);
   U6560 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_5, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_5_port, 
                           B1 => n14, Y => n1808);
   U6561 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn9, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn10, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_5_port);
   U6562 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_8, 
                           B0 => n1806, Y => n1824);
   U6563 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_7, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_7_port, 
                           B1 => n14, Y => n1806);
   U6564 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn5, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn6, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_7_port);
   U6565 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_10, 
                           B0 => n1804, Y => n1822);
   U6566 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_9, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_9_port, 
                           B1 => n14, Y => n1804);
   U6567 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn1, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn2, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_9_port);
   U6568 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_12, 
                           B0 => n1802, Y => n1820);
   U6569 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_11, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_11_port, 
                           B1 => n14, Y => n1802);
   U6570 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn33, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn34, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_11_port);
   U6571 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_14, 
                           B0 => n1800, Y => n1818);
   U6572 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_13, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_13_port, 
                           B1 => n14, Y => n1800);
   U6573 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn29, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn30, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_13_port);
   U6574 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_16, 
                           B0 => n1798, Y => n1816);
   U6575 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_15, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_15_port, 
                           B1 => n14, Y => n1798);
   U6576 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn25, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn26, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_15_port);
   U6577 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_4, 
                           B0 => n1920, Y => n1938);
   U6578 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_3, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_3_port, 
                           B1 => n15, Y => n1920);
   U6579 : XOR2X1 port map( A => n1645, B => n1646, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_3_port);
   U6580 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_6, 
                           B0 => n1918, Y => n1936);
   U6581 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_5, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_5_port, 
                           B1 => n15, Y => n1918);
   U6582 : XOR2X1 port map( A => n1641, B => n1642, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_5_port);
   U6583 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_8, 
                           B0 => n1916, Y => n1934);
   U6584 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_7, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_7_port, 
                           B1 => n15, Y => n1916);
   U6585 : XOR2X1 port map( A => n1637, B => n1638, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_7_port);
   U6586 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_10, 
                           B0 => n1914, Y => n1932);
   U6587 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_9, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_9_port, 
                           B1 => n15, Y => n1914);
   U6588 : XOR2X1 port map( A => n1633, B => n1634, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_9_port);
   U6589 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_12, 
                           B0 => n1912, Y => n1930);
   U6590 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_11, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_11_port, 
                           B1 => n15, Y => n1912);
   U6591 : XOR2X1 port map( A => n1661, B => n1662, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_11_port);
   U6592 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_14, 
                           B0 => n1910, Y => n1928);
   U6593 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_13, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_13_port, 
                           B1 => n15, Y => n1910);
   U6594 : XOR2X1 port map( A => n1657, B => n1658, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_13_port);
   U6595 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_16, 
                           B0 => n1908, Y => n1926);
   U6596 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_15, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_15_port, 
                           B1 => n15, Y => n1908);
   U6597 : XOR2X1 port map( A => n1653, B => n1654, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_15_port);
   U6598 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_4, 
                           B0 => n2029, Y => n2047);
   U6599 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_3, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_3_port, 
                           B1 => n16, Y => n2029);
   U6600 : XOR2X1 port map( A => n1677, B => n1678, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_3_port);
   U6601 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_6, 
                           B0 => n2027, Y => n2045);
   U6602 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_5, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_5_port, 
                           B1 => n16, Y => n2027);
   U6603 : XOR2X1 port map( A => n1673, B => n1674, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_5_port);
   U6604 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_8, 
                           B0 => n2025, Y => n2043);
   U6605 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_7, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_7_port, 
                           B1 => n16, Y => n2025);
   U6606 : XOR2X1 port map( A => n1669, B => n1670, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_7_port);
   U6607 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_10, 
                           B0 => n2023, Y => n2041);
   U6608 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_9, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_9_port, 
                           B1 => n16, Y => n2023);
   U6609 : XOR2X1 port map( A => n1665, B => n1666, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_9_port);
   U6610 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_12, 
                           B0 => n2021, Y => n2039);
   U6611 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_11, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_11_port, 
                           B1 => n16, Y => n2021);
   U6612 : XOR2X1 port map( A => n1693, B => n1694, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_11_port);
   U6613 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_14, 
                           B0 => n2019, Y => n2037);
   U6614 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_13, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_13_port, 
                           B1 => n16, Y => n2019);
   U6615 : XOR2X1 port map( A => n1689, B => n1690, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_13_port);
   U6616 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_16, 
                           B0 => n2017, Y => n2035);
   U6617 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_15, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_15_port, 
                           B1 => n16, Y => n2017);
   U6618 : XOR2X1 port map( A => n1685, B => n1686, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_15_port);
   U6619 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_4, 
                           B0 => n2139, Y => n2157);
   U6620 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_3, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_3_port, 
                           B1 => n17, Y => n2139);
   U6621 : XOR2X1 port map( A => n1709, B => n1710, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_3_port);
   U6622 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_6, 
                           B0 => n2137, Y => n2155);
   U6623 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_5, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_5_port, 
                           B1 => n17, Y => n2137);
   U6624 : XOR2X1 port map( A => n1705, B => n1706, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_5_port);
   U6625 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_8, 
                           B0 => n2135, Y => n2153);
   U6626 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_7, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_7_port, 
                           B1 => n17, Y => n2135);
   U6627 : XOR2X1 port map( A => n1701, B => n1702, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_7_port);
   U6628 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_10, 
                           B0 => n2133, Y => n2151);
   U6629 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_9, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_9_port, 
                           B1 => n17, Y => n2133);
   U6630 : XOR2X1 port map( A => n1697, B => n1698, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_9_port);
   U6631 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_12, 
                           B0 => n2131, Y => n2149);
   U6632 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_11, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_11_port, 
                           B1 => n17, Y => n2131);
   U6633 : XOR2X1 port map( A => n1725, B => n1726, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_11_port);
   U6634 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_14, 
                           B0 => n2129, Y => n2147);
   U6635 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_13, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_13_port, 
                           B1 => n17, Y => n2129);
   U6636 : XOR2X1 port map( A => n1721, B => n1722, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_13_port);
   U6637 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_16, 
                           B0 => n2127, Y => n2145);
   U6638 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_15, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_15_port, 
                           B1 => n17, Y => n2127);
   U6639 : XOR2X1 port map( A => n1717, B => n1718, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_15_port);
   U6640 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_4, 
                           B0 => n2248, Y => n2266);
   U6641 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_3, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_3_port, 
                           B1 => n18, Y => n2248);
   U6642 : XOR2X1 port map( A => n1741, B => n1742, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_3_port);
   U6643 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_6, 
                           B0 => n2246, Y => n2264);
   U6644 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_5, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_5_port, 
                           B1 => n18, Y => n2246);
   U6645 : XOR2X1 port map( A => n1737, B => n1738, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_5_port);
   U6646 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_8, 
                           B0 => n2244, Y => n2262);
   U6647 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_7, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_7_port, 
                           B1 => n18, Y => n2244);
   U6648 : XOR2X1 port map( A => n1733, B => n1734, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_7_port);
   U6649 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_10, 
                           B0 => n2242, Y => n2260);
   U6650 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_9, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_9_port, 
                           B1 => n18, Y => n2242);
   U6651 : XOR2X1 port map( A => n1729, B => n1730, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_9_port);
   U6652 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_12, 
                           B0 => n2240, Y => n2258);
   U6653 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_11, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_11_port, 
                           B1 => n18, Y => n2240);
   U6654 : XOR2X1 port map( A => n1757, B => n1758, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_11_port);
   U6655 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_14, 
                           B0 => n2238, Y => n2256);
   U6656 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_13, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_13_port, 
                           B1 => n18, Y => n2238);
   U6657 : XOR2X1 port map( A => n1753, B => n1754, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_13_port);
   U6658 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_16, 
                           B0 => n2236, Y => n2254);
   U6659 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_15, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_15_port, 
                           B1 => n18, Y => n2236);
   U6660 : XOR2X1 port map( A => n1749, B => n1750, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_15_port);
   U6661 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_2, 
                           B0 => n1812, Y => n1830);
   U6662 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_1, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_1_port, 
                           B1 => n14, Y => n1812);
   U6663 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn17, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn18, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_1_port);
   U6664 : AND2X2 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_0, B 
                           => n846, Y => 
                           input_times_b0_div_componentxUDxactually_substractsxn17);
   U6665 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_2, 
                           B0 => n1922, Y => n1940);
   U6666 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_1, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_1_port, 
                           B1 => n15, Y => n1922);
   U6667 : XOR2X1 port map( A => n1649, B => n1650, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_1_port);
   U6668 : AND2X2 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_0, B 
                           => n1005, Y => n1649);
   U6669 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_2, 
                           B0 => n2031, Y => n2049);
   U6670 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_1, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_1_port, 
                           B1 => n16, Y => n2031);
   U6671 : XOR2X1 port map( A => n1681, B => n1682, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_1_port);
   U6672 : AND2X2 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_0, B 
                           => n1164, Y => n1681);
   U6673 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_2, 
                           B0 => n2141, Y => n2159);
   U6674 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_1, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_1_port, 
                           B1 => n17, Y => n2141);
   U6675 : XOR2X1 port map( A => n1713, B => n1714, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_1_port);
   U6676 : AND2X2 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_0, B 
                           => n528, Y => n1713);
   U6677 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_2, 
                           B0 => n2250, Y => n2268);
   U6678 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_1, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_1_port, 
                           B1 => n18, Y => n2250);
   U6679 : XOR2X1 port map( A => n1745, B => n1746, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_1_port);
   U6680 : AND2X2 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_0, B 
                           => n687, Y => n1745);
   U6681 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_1, 
                           B0 => n1813, Y => n1831);
   U6682 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_0, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_0_port, 
                           B1 => n14, Y => n1813);
   U6683 : XOR2X1 port map( A => n846, B => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_0, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_0_port);
   U6684 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_1, 
                           B0 => n1923, Y => n1941);
   U6685 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_0, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_0_port, 
                           B1 => n15, Y => n1923);
   U6686 : XOR2X1 port map( A => n1005, B => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_0, Y 
                           => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_0_port);
   U6687 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_1, 
                           B0 => n2032, Y => n2050);
   U6688 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_0, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_0_port, 
                           B1 => n16, Y => n2032);
   U6689 : XOR2X1 port map( A => n1164, B => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_0, Y 
                           => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_0_port);
   U6690 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_1, 
                           B0 => n2142, Y => n2160);
   U6691 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_0, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_0_port, 
                           B1 => n17, Y => n2142);
   U6692 : XOR2X1 port map( A => n528, B => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_0, Y 
                           => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_0_port);
   U6693 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_1, 
                           B0 => n2251, Y => n2269);
   U6694 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_0, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_0_port, 
                           B1 => n18, Y => n2251);
   U6695 : XOR2X1 port map( A => n687, B => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_0, Y 
                           => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_0_port);
   U6696 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n1811, Y => n1829);
   U6697 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_2_port, 
                           B1 => n14, Y => n1811);
   U6698 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn15, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn16, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_2_port);
   U6699 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n1809, Y => n1827);
   U6700 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_4_port, 
                           B1 => n14, Y => n1809);
   U6701 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn11, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn12, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_4_port);
   U6702 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n1807, Y => n1825);
   U6703 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_6_port, 
                           B1 => n14, Y => n1807);
   U6704 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn7, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn8, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_6_port);
   U6705 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n1805, Y => n1823);
   U6706 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_8_port, 
                           B1 => n14, Y => n1805);
   U6707 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn3, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn4, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_8_port);
   U6708 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n1803, Y => n1821);
   U6709 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_10_port, 
                           B1 => n14, Y => n1803);
   U6710 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn36, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn35, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_10_port);
   U6711 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n1801, Y => n1819);
   U6712 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_12_port, 
                           B1 => n14, Y => n1801);
   U6713 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn32, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn31, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_12_port);
   U6714 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n1799, Y => n1817);
   U6715 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_14_port, 
                           B1 => n14, Y => n1799);
   U6716 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn28, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn27, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_14_port);
   U6717 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n1921, Y => n1939);
   U6718 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_2_port, 
                           B1 => n15, Y => n1921);
   U6719 : XOR2X1 port map( A => n1647, B => n1648, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_2_port);
   U6720 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n1919, Y => n1937);
   U6721 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_4_port, 
                           B1 => n15, Y => n1919);
   U6722 : XOR2X1 port map( A => n1643, B => n1644, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_4_port);
   U6723 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n1917, Y => n1935);
   U6724 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_6_port, 
                           B1 => n15, Y => n1917);
   U6725 : XOR2X1 port map( A => n1639, B => n1640, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_6_port);
   U6726 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n1915, Y => n1933);
   U6727 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_8_port, 
                           B1 => n15, Y => n1915);
   U6728 : XOR2X1 port map( A => n1635, B => n1636, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_8_port);
   U6729 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n1913, Y => n1931);
   U6730 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_10_port, 
                           B1 => n15, Y => n1913);
   U6731 : XOR2X1 port map( A => n1664, B => n1663, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_10_port);
   U6732 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n1911, Y => n1929);
   U6733 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_12_port, 
                           B1 => n15, Y => n1911);
   U6734 : XOR2X1 port map( A => n1660, B => n1659, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_12_port);
   U6735 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n1909, Y => n1927);
   U6736 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_14_port, 
                           B1 => n15, Y => n1909);
   U6737 : XOR2X1 port map( A => n1656, B => n1655, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_14_port);
   U6738 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n2030, Y => n2048);
   U6739 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_2_port, 
                           B1 => n16, Y => n2030);
   U6740 : XOR2X1 port map( A => n1679, B => n1680, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_2_port);
   U6741 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n2028, Y => n2046);
   U6742 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_4_port, 
                           B1 => n16, Y => n2028);
   U6743 : XOR2X1 port map( A => n1675, B => n1676, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_4_port);
   U6744 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n2026, Y => n2044);
   U6745 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_6_port, 
                           B1 => n16, Y => n2026);
   U6746 : XOR2X1 port map( A => n1671, B => n1672, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_6_port);
   U6747 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n2024, Y => n2042);
   U6748 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_8_port, 
                           B1 => n16, Y => n2024);
   U6749 : XOR2X1 port map( A => n1667, B => n1668, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_8_port);
   U6750 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n2022, Y => n2040);
   U6751 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_10_port, 
                           B1 => n16, Y => n2022);
   U6752 : XOR2X1 port map( A => n1696, B => n1695, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_10_port);
   U6753 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n2020, Y => n2038);
   U6754 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_12_port, 
                           B1 => n16, Y => n2020);
   U6755 : XOR2X1 port map( A => n1692, B => n1691, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_12_port);
   U6756 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n2018, Y => n2036);
   U6757 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_14_port, 
                           B1 => n16, Y => n2018);
   U6758 : XOR2X1 port map( A => n1688, B => n1687, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_14_port);
   U6759 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n2140, Y => n2158);
   U6760 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_2_port, 
                           B1 => n17, Y => n2140);
   U6761 : XOR2X1 port map( A => n1711, B => n1712, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_2_port);
   U6762 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n2138, Y => n2156);
   U6763 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_4_port, 
                           B1 => n17, Y => n2138);
   U6764 : XOR2X1 port map( A => n1707, B => n1708, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_4_port);
   U6765 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n2136, Y => n2154);
   U6766 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_6_port, 
                           B1 => n17, Y => n2136);
   U6767 : XOR2X1 port map( A => n1703, B => n1704, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_6_port);
   U6768 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n2134, Y => n2152);
   U6769 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_8_port, 
                           B1 => n17, Y => n2134);
   U6770 : XOR2X1 port map( A => n1699, B => n1700, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_8_port);
   U6771 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n2132, Y => n2150);
   U6772 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_10_port, 
                           B1 => n17, Y => n2132);
   U6773 : XOR2X1 port map( A => n1728, B => n1727, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_10_port);
   U6774 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n2130, Y => n2148);
   U6775 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_12_port, 
                           B1 => n17, Y => n2130);
   U6776 : XOR2X1 port map( A => n1724, B => n1723, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_12_port);
   U6777 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n2128, Y => n2146);
   U6778 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_14_port, 
                           B1 => n17, Y => n2128);
   U6779 : XOR2X1 port map( A => n1720, B => n1719, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_14_port);
   U6780 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_3, 
                           B0 => n2249, Y => n2267);
   U6781 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_2, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_2_port, 
                           B1 => n18, Y => n2249);
   U6782 : XOR2X1 port map( A => n1743, B => n1744, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_2_port);
   U6783 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_5, 
                           B0 => n2247, Y => n2265);
   U6784 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_4, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_4_port, 
                           B1 => n18, Y => n2247);
   U6785 : XOR2X1 port map( A => n1739, B => n1740, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_4_port);
   U6786 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_7, 
                           B0 => n2245, Y => n2263);
   U6787 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_6, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_6_port, 
                           B1 => n18, Y => n2245);
   U6788 : XOR2X1 port map( A => n1735, B => n1736, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_6_port);
   U6789 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_9, 
                           B0 => n2243, Y => n2261);
   U6790 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_8, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_8_port, 
                           B1 => n18, Y => n2243);
   U6791 : XOR2X1 port map( A => n1731, B => n1732, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_8_port);
   U6792 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_11, 
                           B0 => n2241, Y => n2259);
   U6793 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_10, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_10_port, 
                           B1 => n18, Y => n2241);
   U6794 : XOR2X1 port map( A => n1760, B => n1759, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_10_port);
   U6795 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_13, 
                           B0 => n2239, Y => n2257);
   U6796 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_12, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_12_port, 
                           B1 => n18, Y => n2239);
   U6797 : XOR2X1 port map( A => n1756, B => n1755, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_12_port);
   U6798 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_15, 
                           B0 => n2237, Y => n2255);
   U6799 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_14, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_14_port, 
                           B1 => n18, Y => n2237);
   U6800 : XOR2X1 port map( A => n1752, B => n1751, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_14_port);
   U6801 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_0, 
                           B0 => n1814, Y => n1832);
   U6802 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxshifted_substraction_result_0, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxshifted_substraction_result_0, 
                           B1 => n14, Y => n1814);
   U6803 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_0, 
                           B0 => n1924, Y => n1942);
   U6804 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxshifted_substraction_result_0, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxshifted_substraction_result_0, 
                           B1 => n15, Y => n1924);
   U6805 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_0, 
                           B0 => n2033, Y => n2051);
   U6806 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxshifted_substraction_result_0, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxshifted_substraction_result_0, 
                           B1 => n16, Y => n2033);
   U6807 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_0, 
                           B0 => n2143, Y => n2161);
   U6808 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxshifted_substraction_result_0, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxshifted_substraction_result_0, 
                           B1 => n17, Y => n2143);
   U6809 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_0, 
                           B0 => n2252, Y => n2270);
   U6810 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxshifted_substraction_result_0, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxshifted_substraction_result_0, 
                           B1 => n18, Y => n2252);
   U6811 : OAI2BB1X1 port map( A0N => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_17, 
                           A1N => n371, B0 => n1797, Y => n1815);
   U6812 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_16, 
                           A1 => n2, B0 => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_16_port, 
                           B1 => n14, Y => n1797);
   U6813 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxactually_substractsxn24, B 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn23, Y 
                           => 
                           input_times_b0_div_componentxUDxsubstraction_result_too_long_16_port);
   U6814 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_16, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_16_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn24);
   U6815 : OAI2BB1X1 port map( A0N => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_17, 
                           A1N => n367, B0 => n1907, Y => n1925);
   U6816 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_16, 
                           A1 => n3, B0 => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_16_port, 
                           B1 => n15, Y => n1907);
   U6817 : XOR2X1 port map( A => n1652, B => n1651, Y => 
                           input_p1_times_b1_div_componentxUDxsubstraction_result_too_long_16_port);
   U6818 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_16, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_16_port, Y 
                           => n1652);
   U6819 : OAI2BB1X1 port map( A0N => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_17, 
                           A1N => n372, B0 => n2016, Y => n2034);
   U6820 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_16, 
                           A1 => n4, B0 => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_16_port, 
                           B1 => n16, Y => n2016);
   U6821 : XOR2X1 port map( A => n1684, B => n1683, Y => 
                           input_p2_times_b2_div_componentxUDxsubstraction_result_too_long_16_port);
   U6822 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_16, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_16_port, Y 
                           => n1684);
   U6823 : OAI2BB1X1 port map( A0N => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_17, 
                           A1N => n370, B0 => n2126, Y => n2144);
   U6824 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_16, 
                           A1 => n5, B0 => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_16_port, 
                           B1 => n17, Y => n2126);
   U6825 : XOR2X1 port map( A => n1716, B => n1715, Y => 
                           output_p1_times_a1_div_componentxUDxsubstraction_result_too_long_16_port);
   U6826 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_16, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_16_port, Y 
                           => n1716);
   U6827 : OAI2BB1X1 port map( A0N => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_17, 
                           A1N => n367, B0 => n2235, Y => n2253);
   U6828 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_16, 
                           A1 => n6, B0 => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_16_port, 
                           B1 => n18, Y => n2235);
   U6829 : XOR2X1 port map( A => n1748, B => n1747, Y => 
                           output_p2_times_a2_div_componentxUDxsubstraction_result_too_long_16_port);
   U6830 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_16, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_16_port, Y 
                           => n1748);
   U6831 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_5, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_5_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn10);
   U6832 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_5, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_5_port, Y 
                           => n1642);
   U6833 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_5, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_5_port, Y 
                           => n1674);
   U6834 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_5, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_5_port, Y 
                           => n1706);
   U6835 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_5, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_5_port, Y 
                           => n1738);
   U6836 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_7, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_7_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn6);
   U6837 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_7, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_7_port, Y 
                           => n1638);
   U6838 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_7, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_7_port, Y 
                           => n1670);
   U6839 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_7, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_7_port, Y 
                           => n1702);
   U6840 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_7, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_7_port, Y 
                           => n1734);
   U6841 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_4, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_4_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn11);
   U6842 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_4, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_4_port, Y 
                           => n1643);
   U6843 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_4, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_4_port, Y 
                           => n1675);
   U6844 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_4, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_4_port, Y 
                           => n1707);
   U6845 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_4, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_4_port, Y 
                           => n1739);
   U6846 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_6, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_6_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn7);
   U6847 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_6, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_6_port, Y 
                           => n1639);
   U6848 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_6, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_6_port, Y 
                           => n1671);
   U6849 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_6, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_6_port, Y 
                           => n1703);
   U6850 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_6, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_6_port, Y 
                           => n1735);
   U6851 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_0_port, 
                           B0 => n1850, Y => n1868);
   U6852 : NAND2X1 port map( A => n837, B => en, Y => n1850);
   U6853 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_0_port, 
                           B0 => n1960, Y => n1978);
   U6854 : NAND2X1 port map( A => n996, B => en, Y => n1960);
   U6855 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_0_port, 
                           B0 => n2069, Y => n2087);
   U6856 : NAND2X1 port map( A => n1155, B => en, Y => n2069);
   U6857 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_0_port, 
                           B0 => n2179, Y => n2197);
   U6858 : NAND2X1 port map( A => n519, B => en, Y => n2179);
   U6859 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_0_port, 
                           B0 => n2288, Y => n2306);
   U6860 : NAND2X1 port map( A => n678, B => en, Y => n2288);
   U6861 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_9, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_9_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn2);
   U6862 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_9, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_9_port, Y 
                           => n1634);
   U6863 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_9, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_9_port, Y 
                           => n1666);
   U6864 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_9, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_9_port, Y 
                           => n1698);
   U6865 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_9, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_9_port, Y 
                           => n1730);
   U6866 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_11, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_11_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn34);
   U6867 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_11, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_11_port, Y 
                           => n1662);
   U6868 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_11, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_11_port, Y 
                           => n1694);
   U6869 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_11, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_11_port, Y 
                           => n1726);
   U6870 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_11, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_11_port, Y 
                           => n1758);
   U6871 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_8, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_8_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn3);
   U6872 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_8, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_8_port, Y 
                           => n1635);
   U6873 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_8, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_8_port, Y 
                           => n1667);
   U6874 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_8, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_8_port, Y 
                           => n1699);
   U6875 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_8, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_8_port, Y 
                           => n1731);
   U6876 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_10, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_10_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn36);
   U6877 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_10, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_10_port, Y 
                           => n1664);
   U6878 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_10, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_10_port, Y 
                           => n1696);
   U6879 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_10, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_10_port, Y 
                           => n1728);
   U6880 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_10, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_10_port, Y 
                           => n1760);
   U6881 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_12, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_12_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn32);
   U6882 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_12, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_12_port, Y 
                           => n1660);
   U6883 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_12, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_12_port, Y 
                           => n1692);
   U6884 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_12, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_12_port, Y 
                           => n1724);
   U6885 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_12, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_12_port, Y 
                           => n1756);
   U6886 : INVX1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_9, Y 
                           => n1529);
   U6887 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_9, Y 
                           => n1513);
   U6888 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_9, Y 
                           => n1497);
   U6889 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_9, Y 
                           => n1481);
   U6890 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_9, Y 
                           => n1465);
   U6891 : BUFX4 port map( A => n4673, Y => change_input_port);
   U6892 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_13, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_13_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn30);
   U6893 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_13, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_13_port, Y 
                           => n1658);
   U6894 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_13, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_13_port, Y 
                           => n1690);
   U6895 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_13, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_13_port, Y 
                           => n1722);
   U6896 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_13, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_13_port, Y 
                           => n1754);
   U6897 : XOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_15, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_15_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn26);
   U6898 : XOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_15, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_15_port, Y 
                           => n1654);
   U6899 : XOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_15, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_15_port, Y 
                           => n1686);
   U6900 : XOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_15, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_15_port, Y 
                           => n1718);
   U6901 : XOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_15, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_15_port, Y 
                           => n1750);
   U6902 : XNOR2X1 port map( A => 
                           input_times_b0_div_componentxUDxcentral_parallel_output_14, B 
                           => 
                           input_times_b0_div_componentxUDxsub_ready_negative_divisor_14_port, Y 
                           => 
                           input_times_b0_div_componentxUDxactually_substractsxn28);
   U6903 : XNOR2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxcentral_parallel_output_14, B 
                           => 
                           input_p1_times_b1_div_componentxUDxsub_ready_negative_divisor_14_port, Y 
                           => n1656);
   U6904 : XNOR2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxcentral_parallel_output_14, B 
                           => 
                           input_p2_times_b2_div_componentxUDxsub_ready_negative_divisor_14_port, Y 
                           => n1688);
   U6905 : XNOR2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxcentral_parallel_output_14, B 
                           => 
                           output_p1_times_a1_div_componentxUDxsub_ready_negative_divisor_14_port, Y 
                           => n1720);
   U6906 : XNOR2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxcentral_parallel_output_14, B 
                           => 
                           output_p2_times_a2_div_componentxUDxsub_ready_negative_divisor_14_port, Y 
                           => n1752);
   U6907 : OAI2BB2X1 port map( B0 => n1191, B1 => n321, A0N => 
                           input_previous_1_9_port, A1N => n321, Y => n4628);
   U6908 : OAI2BB2X1 port map( B0 => n1293, B1 => n1260, A0N => 
                           input_previous_2_9_port, A1N => n320, Y => n4646);
   U6909 : OAI2BB2X1 port map( B0 => n1198, B1 => n1260, A0N => 
                           input_previous_1_16_port, A1N => n321, Y => n4635);
   U6910 : INVX1 port map( A => input_previous_0_16_port, Y => n1198);
   U6911 : OAI2BB2X1 port map( B0 => n1197, B1 => n1260, A0N => 
                           input_previous_1_15_port, A1N => n321, Y => n4634);
   U6912 : INVX1 port map( A => input_previous_0_15_port, Y => n1197);
   U6913 : OAI2BB2X1 port map( B0 => n1196, B1 => n320, A0N => 
                           input_previous_1_14_port, A1N => n321, Y => n4633);
   U6914 : INVX1 port map( A => input_previous_0_14_port, Y => n1196);
   U6915 : OAI2BB2X1 port map( B0 => n1195, B1 => n1260, A0N => 
                           input_previous_1_13_port, A1N => n321, Y => n4632);
   U6916 : INVX1 port map( A => input_previous_0_13_port, Y => n1195);
   U6917 : OAI2BB2X1 port map( B0 => n1194, B1 => n1260, A0N => 
                           input_previous_1_12_port, A1N => n321, Y => n4631);
   U6918 : INVX1 port map( A => input_previous_0_12_port, Y => n1194);
   U6919 : OAI2BB2X1 port map( B0 => n1193, B1 => n319, A0N => 
                           input_previous_1_11_port, A1N => n321, Y => n4630);
   U6920 : INVX1 port map( A => input_previous_0_11_port, Y => n1193);
   U6921 : OAI2BB2X1 port map( B0 => n1192, B1 => n319, A0N => 
                           input_previous_1_10_port, A1N => n321, Y => n4629);
   U6922 : INVX1 port map( A => input_previous_0_10_port, Y => n1192);
   U6923 : OAI2BB2X1 port map( B0 => n1190, B1 => n1260, A0N => 
                           input_previous_1_8_port, A1N => n321, Y => n4627);
   U6924 : INVX1 port map( A => input_previous_0_8_port, Y => n1190);
   U6925 : OAI2BB2X1 port map( B0 => n1189, B1 => n1260, A0N => 
                           input_previous_1_7_port, A1N => n321, Y => n4626);
   U6926 : INVX1 port map( A => input_previous_0_7_port, Y => n1189);
   U6927 : OAI2BB2X1 port map( B0 => n1188, B1 => n1260, A0N => 
                           input_previous_1_6_port, A1N => n321, Y => n4625);
   U6928 : INVX1 port map( A => input_previous_0_6_port, Y => n1188);
   U6929 : OAI2BB2X1 port map( B0 => n1187, B1 => n321, A0N => 
                           input_previous_1_5_port, A1N => n321, Y => n4624);
   U6930 : INVX1 port map( A => input_previous_0_5_port, Y => n1187);
   U6931 : OAI2BB2X1 port map( B0 => n1186, B1 => n1260, A0N => 
                           input_previous_1_4_port, A1N => n321, Y => n4623);
   U6932 : INVX1 port map( A => input_previous_0_4_port, Y => n1186);
   U6933 : OAI2BB2X1 port map( B0 => n1185, B1 => n1260, A0N => 
                           input_previous_1_3_port, A1N => n321, Y => n4622);
   U6934 : INVX1 port map( A => input_previous_0_3_port, Y => n1185);
   U6935 : OAI2BB2X1 port map( B0 => n1184, B1 => n1260, A0N => 
                           input_previous_1_2_port, A1N => n321, Y => n4621);
   U6936 : INVX1 port map( A => input_previous_0_2_port, Y => n1184);
   U6937 : OAI2BB2X1 port map( B0 => n1183, B1 => n321, A0N => 
                           input_previous_1_1_port, A1N => n321, Y => n4620);
   U6938 : INVX1 port map( A => input_previous_0_1_port, Y => n1183);
   U6939 : OAI2BB2X1 port map( B0 => n1182, B1 => n1260, A0N => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_0_port, 
                           A1N => n319, Y => n4619);
   U6940 : INVX1 port map( A => 
                           input_times_b0_mul_componentxinput_A_inverted_0_port
                           , Y => n1182);
   U6941 : OAI2BB2X1 port map( B0 => n1300, B1 => n1260, A0N => 
                           input_previous_2_16_port, A1N => n320, Y => n4653);
   U6942 : INVX1 port map( A => input_previous_1_16_port, Y => n1300);
   U6943 : OAI2BB2X1 port map( B0 => n1299, B1 => n1260, A0N => 
                           input_previous_2_15_port, A1N => n320, Y => n4652);
   U6944 : INVX1 port map( A => input_previous_1_15_port, Y => n1299);
   U6945 : OAI2BB2X1 port map( B0 => n1298, B1 => n1260, A0N => 
                           input_previous_2_14_port, A1N => n320, Y => n4651);
   U6946 : INVX1 port map( A => input_previous_1_14_port, Y => n1298);
   U6947 : OAI2BB2X1 port map( B0 => n1297, B1 => n321, A0N => 
                           input_previous_2_13_port, A1N => n320, Y => n4650);
   U6948 : INVX1 port map( A => input_previous_1_13_port, Y => n1297);
   U6949 : OAI2BB2X1 port map( B0 => n1296, B1 => n1260, A0N => 
                           input_previous_2_12_port, A1N => n320, Y => n4649);
   U6950 : INVX1 port map( A => input_previous_1_12_port, Y => n1296);
   U6951 : OAI2BB2X1 port map( B0 => n1295, B1 => n1260, A0N => 
                           input_previous_2_11_port, A1N => n320, Y => n4648);
   U6952 : INVX1 port map( A => input_previous_1_11_port, Y => n1295);
   U6953 : OAI2BB2X1 port map( B0 => n1294, B1 => n320, A0N => 
                           input_previous_2_10_port, A1N => n320, Y => n4647);
   U6954 : INVX1 port map( A => input_previous_1_10_port, Y => n1294);
   U6955 : OAI2BB2X1 port map( B0 => n1292, B1 => n1260, A0N => 
                           input_previous_2_8_port, A1N => n320, Y => n4645);
   U6956 : INVX1 port map( A => input_previous_1_8_port, Y => n1292);
   U6957 : OAI2BB2X1 port map( B0 => n1291, B1 => n319, A0N => 
                           input_previous_2_7_port, A1N => n320, Y => n4644);
   U6958 : INVX1 port map( A => input_previous_1_7_port, Y => n1291);
   U6959 : OAI2BB2X1 port map( B0 => n1290, B1 => n321, A0N => 
                           input_previous_2_6_port, A1N => n321, Y => n4643);
   U6960 : INVX1 port map( A => input_previous_1_6_port, Y => n1290);
   U6961 : OAI2BB2X1 port map( B0 => n1289, B1 => n320, A0N => 
                           input_previous_2_5_port, A1N => n321, Y => n4642);
   U6962 : INVX1 port map( A => input_previous_1_5_port, Y => n1289);
   U6963 : OAI2BB2X1 port map( B0 => n1288, B1 => n319, A0N => 
                           input_previous_2_4_port, A1N => n321, Y => n4641);
   U6964 : INVX1 port map( A => input_previous_1_4_port, Y => n1288);
   U6965 : OAI2BB2X1 port map( B0 => n1287, B1 => n321, A0N => 
                           input_previous_2_3_port, A1N => n321, Y => n4640);
   U6966 : INVX1 port map( A => input_previous_1_3_port, Y => n1287);
   U6967 : OAI2BB2X1 port map( B0 => n1286, B1 => n320, A0N => 
                           input_previous_2_2_port, A1N => n321, Y => n4639);
   U6968 : INVX1 port map( A => input_previous_1_2_port, Y => n1286);
   U6969 : OAI2BB2X1 port map( B0 => n1285, B1 => n320, A0N => 
                           input_previous_2_1_port, A1N => n321, Y => n4638);
   U6970 : INVX1 port map( A => input_previous_1_1_port, Y => n1285);
   U6971 : OAI2BB2X1 port map( B0 => n1284, B1 => n319, A0N => 
                           input_p2_times_b2_mul_componentxinput_A_inverted_0_port, 
                           A1N => n321, Y => n4637);
   U6972 : INVX1 port map( A => 
                           input_p1_times_b1_mul_componentxinput_A_inverted_0_port, Y 
                           => n1284);
   U6973 : OAI2BB2X1 port map( B0 => n1174, B1 => n320, A0N => 
                           input_previous_0_16_port, A1N => n319, Y => 
                           input_prev_0_registerxn18);
   U6974 : OAI2BB2X1 port map( B0 => n1174, B1 => n321, A0N => 
                           input_previous_0_15_port, A1N => n320, Y => 
                           input_prev_0_registerxn17);
   U6975 : OAI2BB2X1 port map( B0 => n1174, B1 => n1260, A0N => 
                           input_previous_0_14_port, A1N => n319, Y => 
                           input_prev_0_registerxn16);
   U6976 : OAI2BB2X1 port map( B0 => n1174, B1 => n321, A0N => 
                           input_previous_0_13_port, A1N => n319, Y => 
                           input_prev_0_registerxn15);
   U6977 : OAI2BB2X1 port map( B0 => n1174, B1 => n1260, A0N => 
                           input_previous_0_12_port, A1N => n319, Y => 
                           input_prev_0_registerxn14);
   U6978 : OAI2BB2X1 port map( B0 => n1174, B1 => n1260, A0N => 
                           input_previous_0_11_port, A1N => n319, Y => 
                           input_prev_0_registerxn13);
   U6979 : OAI2BB2X1 port map( B0 => n1174, B1 => n320, A0N => 
                           input_previous_0_10_port, A1N => n319, Y => 
                           input_prev_0_registerxn12);
   U6980 : OAI2BB2X1 port map( B0 => n1174, B1 => n1260, A0N => 
                           input_previous_0_9_port, A1N => n319, Y => 
                           input_prev_0_registerxn11);
   U6981 : OAI2BB2X1 port map( B0 => n1174, B1 => n321, A0N => 
                           input_previous_0_8_port, A1N => n319, Y => 
                           input_prev_0_registerxn10);
   U6982 : OAI2BB2X1 port map( B0 => n1174, B1 => n320, A0N => 
                           input_previous_0_7_port, A1N => n319, Y => 
                           input_prev_0_registerxn9);
   U6983 : OAI2BB2X1 port map( B0 => n1175, B1 => n319, A0N => 
                           input_previous_0_6_port, A1N => n319, Y => 
                           input_prev_0_registerxn8);
   U6984 : INVX1 port map( A => input_signal(6), Y => n1175);
   U6985 : OAI2BB2X1 port map( B0 => n1176, B1 => n1260, A0N => 
                           input_previous_0_5_port, A1N => n319, Y => 
                           input_prev_0_registerxn7);
   U6986 : INVX1 port map( A => input_signal(5), Y => n1176);
   U6987 : OAI2BB2X1 port map( B0 => n1177, B1 => n1260, A0N => 
                           input_previous_0_4_port, A1N => n319, Y => 
                           input_prev_0_registerxn6);
   U6988 : INVX1 port map( A => input_signal(4), Y => n1177);
   U6989 : OAI2BB2X1 port map( B0 => n1178, B1 => n321, A0N => 
                           input_previous_0_3_port, A1N => n319, Y => 
                           input_prev_0_registerxn5);
   U6990 : INVX1 port map( A => input_signal(3), Y => n1178);
   U6991 : OAI2BB2X1 port map( B0 => n1179, B1 => n1260, A0N => 
                           input_previous_0_2_port, A1N => n319, Y => 
                           input_prev_0_registerxn4);
   U6992 : INVX1 port map( A => input_signal(2), Y => n1179);
   U6993 : OAI2BB2X1 port map( B0 => n1180, B1 => n319, A0N => 
                           input_previous_0_1_port, A1N => n319, Y => 
                           input_prev_0_registerxn3);
   U6994 : INVX1 port map( A => input_signal(1), Y => n1180);
   U6995 : OAI2BB2X1 port map( B0 => n1181, B1 => n1260, A0N => 
                           input_times_b0_mul_componentxinput_A_inverted_0_port
                           , A1N => n319, Y => input_prev_0_registerxn2);
   U6996 : INVX1 port map( A => input_signal(0), Y => n1181);
   U6997 : NAND2X1 port map( A => change_input_port, B => en, Y => n109);
   U6998 : INVX1 port map( A => n109, Y => n1871);
   U6999 : NAND2X1 port map( A => change_input_port, B => en, Y => n110);
   U7000 : INVX1 port map( A => n110, Y => n2090);
   U7001 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           B => en, Y => n4203);
   U7002 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           B => en, Y => n4259);
   U7003 : NAND2X1 port map( A => n7, B => en, Y => n4369);
   U7004 : NAND2X1 port map( A => n8, B => en, Y => 
                           input_times_b0_div_componentxn24);
   U7005 : OAI22X1 port map( A0 => n374, A1 => n151, B0 => n1381, B1 => n4203, 
                           Y => n4240);
   U7006 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxoutput_sign_gated_prev, Y 
                           => n1381);
   U7007 : OAI22X1 port map( A0 => n376, A1 => n149, B0 => n1361, B1 => n4259, 
                           Y => n4296);
   U7008 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxoutput_sign_gated_prev, Y 
                           => n1361);
   U7009 : OAI22X1 port map( A0 => n378, A1 => n145, B0 => n1322, B1 => n4369, 
                           Y => n4406);
   U7010 : INVX1 port map( A => 
                           output_p2_times_a2_div_componentxoutput_sign_gated_prev, Y 
                           => n1322);
   U7011 : OAI22X1 port map( A0 => n380, A1 => n135, B0 => n1239, B1 => 
                           input_times_b0_div_componentxn24, Y => 
                           input_times_b0_div_componentxn62);
   U7012 : INVX1 port map( A => 
                           input_times_b0_div_componentxoutput_sign_gated_prev,
                           Y => n1239);
   U7013 : OAI22X1 port map( A0 => n367, A1 => n1252, B0 => en, B1 => n1251, Y 
                           => clock_chopper_and_divisionxn37);
   U7014 : OAI22X1 port map( A0 => en, A1 => n1240, B0 => n1241, B1 => n367, Y 
                           => clock_chopper_and_divisionxn26);
   U7015 : OAI22X1 port map( A0 => en, A1 => n1259, B0 => n367, B1 => n1261, Y 
                           => clock_chopper_and_divisionxn45);
   U7016 : OAI22X1 port map( A0 => en, A1 => n1258, B0 => n368, B1 => n1259, Y 
                           => clock_chopper_and_divisionxn44);
   U7017 : OAI22X1 port map( A0 => en, A1 => n1257, B0 => n367, B1 => n1258, Y 
                           => clock_chopper_and_divisionxn43);
   U7018 : OAI22X1 port map( A0 => en, A1 => n1256, B0 => n367, B1 => n1257, Y 
                           => clock_chopper_and_divisionxn42);
   U7019 : OAI22X1 port map( A0 => en, A1 => n1255, B0 => n367, B1 => n1256, Y 
                           => clock_chopper_and_divisionxn41);
   U7020 : OAI22X1 port map( A0 => en, A1 => n1254, B0 => n370, B1 => n1255, Y 
                           => clock_chopper_and_divisionxn40);
   U7021 : OAI22X1 port map( A0 => en, A1 => n1253, B0 => n367, B1 => n1254, Y 
                           => clock_chopper_and_divisionxn39);
   U7022 : OAI22X1 port map( A0 => en, A1 => n1252, B0 => n369, B1 => n1253, Y 
                           => clock_chopper_and_divisionxn38);
   U7023 : OAI22X1 port map( A0 => en, A1 => n1250, B0 => n368, B1 => n1251, Y 
                           => clock_chopper_and_divisionxn36);
   U7024 : OAI22X1 port map( A0 => en, A1 => n1249, B0 => n367, B1 => n1250, Y 
                           => clock_chopper_and_divisionxn35);
   U7025 : OAI22X1 port map( A0 => en, A1 => n1248, B0 => n369, B1 => n1249, Y 
                           => clock_chopper_and_divisionxn34);
   U7026 : OAI22X1 port map( A0 => en, A1 => n1247, B0 => n368, B1 => n1248, Y 
                           => clock_chopper_and_divisionxn33);
   U7027 : OAI22X1 port map( A0 => en, A1 => n1246, B0 => n367, B1 => n1247, Y 
                           => clock_chopper_and_divisionxn32);
   U7028 : OAI22X1 port map( A0 => en, A1 => n1245, B0 => n367, B1 => n1246, Y 
                           => clock_chopper_and_divisionxn31);
   U7029 : OAI22X1 port map( A0 => en, A1 => n1244, B0 => n367, B1 => n1245, Y 
                           => clock_chopper_and_divisionxn30);
   U7030 : OAI22X1 port map( A0 => en, A1 => n1243, B0 => n367, B1 => n1244, Y 
                           => clock_chopper_and_divisionxn29);
   U7031 : OAI22X1 port map( A0 => en, A1 => n1242, B0 => n367, B1 => n1243, Y 
                           => clock_chopper_and_divisionxn28);
   U7032 : OAI22X1 port map( A0 => en, A1 => n1241, B0 => n367, B1 => n1242, Y 
                           => clock_chopper_and_divisionxn27);
   U7033 : OAI22X1 port map( A0 => n367, A1 => n1240, B0 => en, B1 => n1262, Y 
                           => clock_chopper_and_divisionxn49);
   U7034 : OAI22X1 port map( A0 => en, A1 => n1261, B0 => n367, B1 => n1262, Y 
                           => clock_chopper_and_divisionxn47);
   U7035 : INVX1 port map( A => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n161);
   U7036 : INVX1 port map( A => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n162);
   U7037 : INVX1 port map( A => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n163);
   U7038 : OAI2BB2X1 port map( B0 => n367, B1 => n1261, A0N => n258, A1N => 
                           n368, Y => clock_chopper_and_divisionxn46);
   U7039 : BUFX3 port map( A => n4673, Y => n258);
   U7040 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_20_port, Y 
                           => n1241);
   U7041 : INVX1 port map( A => clock_chopper_and_divisionxdivision_ring_9_port
                           , Y => n1252);
   U7042 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_21_port, Y 
                           => n1240);
   U7043 : INVX1 port map( A => clock_chopper_and_divisionxdivision_ring_2_port
                           , Y => n1259);
   U7044 : INVX1 port map( A => clock_chopper_and_divisionxdivision_ring_3_port
                           , Y => n1258);
   U7045 : INVX1 port map( A => clock_chopper_and_divisionxdivision_ring_4_port
                           , Y => n1257);
   U7046 : INVX1 port map( A => clock_chopper_and_divisionxdivision_ring_5_port
                           , Y => n1256);
   U7047 : INVX1 port map( A => clock_chopper_and_divisionxdivision_ring_6_port
                           , Y => n1255);
   U7048 : INVX1 port map( A => clock_chopper_and_divisionxdivision_ring_7_port
                           , Y => n1254);
   U7049 : INVX1 port map( A => clock_chopper_and_divisionxdivision_ring_8_port
                           , Y => n1253);
   U7050 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_11_port, Y 
                           => n1250);
   U7051 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_12_port, Y 
                           => n1249);
   U7052 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_13_port, Y 
                           => n1248);
   U7053 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_14_port, Y 
                           => n1247);
   U7054 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_15_port, Y 
                           => n1246);
   U7055 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_16_port, Y 
                           => n1245);
   U7056 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_17_port, Y 
                           => n1244);
   U7057 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_18_port, Y 
                           => n1243);
   U7058 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_19_port, Y 
                           => n1242);
   U7059 : INVX1 port map( A => 
                           clock_chopper_and_divisionxdivision_ring_10_port, Y 
                           => n1251);
   U7060 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_1_port, 
                           B0 => n1849, Y => n1867);
   U7061 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_0_port, B 
                           => en, Y => n1849);
   U7062 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_2_port, 
                           B0 => n1848, Y => n1866);
   U7063 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_1_port, B 
                           => en, Y => n1848);
   U7064 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_3_port, 
                           B0 => n1847, Y => n1865);
   U7065 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_2_port, B 
                           => en, Y => n1847);
   U7066 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_4_port, 
                           B0 => n1846, Y => n1864);
   U7067 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_3_port, B 
                           => en, Y => n1846);
   U7068 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_5_port, 
                           B0 => n1845, Y => n1863);
   U7069 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_4_port, B 
                           => en, Y => n1845);
   U7070 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_6_port, 
                           B0 => n1844, Y => n1862);
   U7071 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_5_port, B 
                           => en, Y => n1844);
   U7072 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_7_port, 
                           B0 => n1843, Y => n1861);
   U7073 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_6_port, B 
                           => en, Y => n1843);
   U7074 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_8_port, 
                           B0 => n1842, Y => n1860);
   U7075 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_7_port, B 
                           => en, Y => n1842);
   U7076 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_9_port, 
                           B0 => n1841, Y => n1859);
   U7077 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_8_port, B 
                           => en, Y => n1841);
   U7078 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_10_port, 
                           B0 => n1840, Y => n1858);
   U7079 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_9_port, B 
                           => en, Y => n1840);
   U7080 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_11_port, 
                           B0 => n1839, Y => n1857);
   U7081 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_10_port, B 
                           => en, Y => n1839);
   U7082 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_12_port, 
                           B0 => n1838, Y => n1856);
   U7083 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_11_port, B 
                           => en, Y => n1838);
   U7084 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_13_port, 
                           B0 => n1837, Y => n1855);
   U7085 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_12_port, B 
                           => en, Y => n1837);
   U7086 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_14_port, 
                           B0 => n1836, Y => n1854);
   U7087 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_13_port, B 
                           => en, Y => n1836);
   U7088 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_15_port, 
                           B0 => n1835, Y => n1853);
   U7089 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_14_port, B 
                           => en, Y => n1835);
   U7090 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_16_port, 
                           B0 => n1834, Y => n1852);
   U7091 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_15_port, B 
                           => en, Y => n1834);
   U7092 : OAI2BB1X1 port map( A0N => 
                           input_times_b0_div_componentxUDxquotient_not_gated_17_port, 
                           A1N => n370, B0 => n1833, Y => n1851);
   U7093 : NAND2X1 port map( A => 
                           input_times_b0_div_componentxUDxquotient_not_gated_16_port, B 
                           => en, Y => n1833);
   U7094 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_1_port, 
                           B0 => n1959, Y => n1977);
   U7095 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_0_port, B 
                           => en, Y => n1959);
   U7096 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_2_port, 
                           B0 => n1958, Y => n1976);
   U7097 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_1_port, B 
                           => en, Y => n1958);
   U7098 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_3_port, 
                           B0 => n1957, Y => n1975);
   U7099 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_2_port, B 
                           => en, Y => n1957);
   U7100 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_4_port, 
                           B0 => n1956, Y => n1974);
   U7101 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_3_port, B 
                           => en, Y => n1956);
   U7102 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_5_port, 
                           B0 => n1955, Y => n1973);
   U7103 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_4_port, B 
                           => en, Y => n1955);
   U7104 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_6_port, 
                           B0 => n1954, Y => n1972);
   U7105 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_5_port, B 
                           => en, Y => n1954);
   U7106 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_7_port, 
                           B0 => n1953, Y => n1971);
   U7107 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_6_port, B 
                           => en, Y => n1953);
   U7108 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_8_port, 
                           B0 => n1952, Y => n1970);
   U7109 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_7_port, B 
                           => en, Y => n1952);
   U7110 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_9_port, 
                           B0 => n1951, Y => n1969);
   U7111 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_8_port, B 
                           => en, Y => n1951);
   U7112 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_10_port, 
                           B0 => n1950, Y => n1968);
   U7113 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_9_port, B 
                           => en, Y => n1950);
   U7114 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_11_port, 
                           B0 => n1949, Y => n1967);
   U7115 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_10_port, B 
                           => en, Y => n1949);
   U7116 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_12_port, 
                           B0 => n1948, Y => n1966);
   U7117 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_11_port, B 
                           => en, Y => n1948);
   U7118 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_13_port, 
                           B0 => n1947, Y => n1965);
   U7119 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_12_port, B 
                           => en, Y => n1947);
   U7120 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_14_port, 
                           B0 => n1946, Y => n1964);
   U7121 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_13_port, B 
                           => en, Y => n1946);
   U7122 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_15_port, 
                           B0 => n1945, Y => n1963);
   U7123 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_14_port, B 
                           => en, Y => n1945);
   U7124 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_16_port, 
                           B0 => n1944, Y => n1962);
   U7125 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_15_port, B 
                           => en, Y => n1944);
   U7126 : OAI2BB1X1 port map( A0N => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_17_port, 
                           A1N => n369, B0 => n1943, Y => n1961);
   U7127 : NAND2X1 port map( A => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_16_port, B 
                           => en, Y => n1943);
   U7128 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_1_port, 
                           B0 => n2068, Y => n2086);
   U7129 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_0_port, B 
                           => en, Y => n2068);
   U7130 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_2_port, 
                           B0 => n2067, Y => n2085);
   U7131 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_1_port, B 
                           => en, Y => n2067);
   U7132 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_3_port, 
                           B0 => n2066, Y => n2084);
   U7133 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_2_port, B 
                           => en, Y => n2066);
   U7134 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_4_port, 
                           B0 => n2065, Y => n2083);
   U7135 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_3_port, B 
                           => en, Y => n2065);
   U7136 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_5_port, 
                           B0 => n2064, Y => n2082);
   U7137 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_4_port, B 
                           => en, Y => n2064);
   U7138 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_6_port, 
                           B0 => n2063, Y => n2081);
   U7139 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_5_port, B 
                           => en, Y => n2063);
   U7140 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_7_port, 
                           B0 => n2062, Y => n2080);
   U7141 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_6_port, B 
                           => en, Y => n2062);
   U7142 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_8_port, 
                           B0 => n2061, Y => n2079);
   U7143 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_7_port, B 
                           => en, Y => n2061);
   U7144 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_9_port, 
                           B0 => n2060, Y => n2078);
   U7145 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_8_port, B 
                           => en, Y => n2060);
   U7146 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_10_port, 
                           B0 => n2059, Y => n2077);
   U7147 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_9_port, B 
                           => en, Y => n2059);
   U7148 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_11_port, 
                           B0 => n2058, Y => n2076);
   U7149 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_10_port, B 
                           => en, Y => n2058);
   U7150 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_12_port, 
                           B0 => n2057, Y => n2075);
   U7151 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_11_port, B 
                           => en, Y => n2057);
   U7152 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_13_port, 
                           B0 => n2056, Y => n2074);
   U7153 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_12_port, B 
                           => en, Y => n2056);
   U7154 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_14_port, 
                           B0 => n2055, Y => n2073);
   U7155 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_13_port, B 
                           => en, Y => n2055);
   U7156 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_15_port, 
                           B0 => n2054, Y => n2072);
   U7157 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_14_port, B 
                           => en, Y => n2054);
   U7158 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_16_port, 
                           B0 => n2053, Y => n2071);
   U7159 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_15_port, B 
                           => en, Y => n2053);
   U7160 : OAI2BB1X1 port map( A0N => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_17_port, 
                           A1N => n369, B0 => n2052, Y => n2070);
   U7161 : NAND2X1 port map( A => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_16_port, B 
                           => en, Y => n2052);
   U7162 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_1_port, 
                           B0 => n2178, Y => n2196);
   U7163 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_0_port, B 
                           => en, Y => n2178);
   U7164 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_2_port, 
                           B0 => n2177, Y => n2195);
   U7165 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_1_port, B 
                           => en, Y => n2177);
   U7166 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_3_port, 
                           B0 => n2176, Y => n2194);
   U7167 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_2_port, B 
                           => en, Y => n2176);
   U7168 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_4_port, 
                           B0 => n2175, Y => n2193);
   U7169 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_3_port, B 
                           => en, Y => n2175);
   U7170 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_5_port, 
                           B0 => n2174, Y => n2192);
   U7171 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_4_port, B 
                           => en, Y => n2174);
   U7172 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_6_port, 
                           B0 => n2173, Y => n2191);
   U7173 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_5_port, B 
                           => en, Y => n2173);
   U7174 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_7_port, 
                           B0 => n2172, Y => n2190);
   U7175 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_6_port, B 
                           => en, Y => n2172);
   U7176 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_8_port, 
                           B0 => n2171, Y => n2189);
   U7177 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_7_port, B 
                           => en, Y => n2171);
   U7178 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_9_port, 
                           B0 => n2170, Y => n2188);
   U7179 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_8_port, B 
                           => en, Y => n2170);
   U7180 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_10_port, 
                           B0 => n2169, Y => n2187);
   U7181 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_9_port, B 
                           => en, Y => n2169);
   U7182 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_11_port, 
                           B0 => n2168, Y => n2186);
   U7183 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_10_port, B 
                           => en, Y => n2168);
   U7184 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_12_port, 
                           B0 => n2167, Y => n2185);
   U7185 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_11_port, B 
                           => en, Y => n2167);
   U7186 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_13_port, 
                           B0 => n2166, Y => n2184);
   U7187 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_12_port, B 
                           => en, Y => n2166);
   U7188 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_14_port, 
                           B0 => n2165, Y => n2183);
   U7189 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_13_port, B 
                           => en, Y => n2165);
   U7190 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_15_port, 
                           B0 => n2164, Y => n2182);
   U7191 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_14_port, B 
                           => en, Y => n2164);
   U7192 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_16_port, 
                           B0 => n2163, Y => n2181);
   U7193 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_15_port, B 
                           => en, Y => n2163);
   U7194 : OAI2BB1X1 port map( A0N => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_17_port, 
                           A1N => n368, B0 => n2162, Y => n2180);
   U7195 : NAND2X1 port map( A => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_16_port, B 
                           => en, Y => n2162);
   U7196 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_1_port, 
                           B0 => n2287, Y => n2305);
   U7197 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_0_port, B 
                           => en, Y => n2287);
   U7198 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_2_port, 
                           B0 => n2286, Y => n2304);
   U7199 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_1_port, B 
                           => en, Y => n2286);
   U7200 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_3_port, 
                           B0 => n2285, Y => n2303);
   U7201 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_2_port, B 
                           => en, Y => n2285);
   U7202 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_4_port, 
                           B0 => n2284, Y => n2302);
   U7203 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_3_port, B 
                           => en, Y => n2284);
   U7204 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_5_port, 
                           B0 => n2283, Y => n2301);
   U7205 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_4_port, B 
                           => en, Y => n2283);
   U7206 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_6_port, 
                           B0 => n2282, Y => n2300);
   U7207 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_5_port, B 
                           => en, Y => n2282);
   U7208 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_7_port, 
                           B0 => n2281, Y => n2299);
   U7209 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_6_port, B 
                           => en, Y => n2281);
   U7210 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_8_port, 
                           B0 => n2280, Y => n2298);
   U7211 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_7_port, B 
                           => en, Y => n2280);
   U7212 : OAI2BB1X1 port map( A0N => n370, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_9_port, 
                           B0 => n2279, Y => n2297);
   U7213 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_8_port, B 
                           => en, Y => n2279);
   U7214 : OAI2BB1X1 port map( A0N => n369, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_10_port, 
                           B0 => n2278, Y => n2296);
   U7215 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_9_port, B 
                           => en, Y => n2278);
   U7216 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_11_port, 
                           B0 => n2277, Y => n2295);
   U7217 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_10_port, B 
                           => en, Y => n2277);
   U7218 : OAI2BB1X1 port map( A0N => n367, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_12_port, 
                           B0 => n2276, Y => n2294);
   U7219 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_11_port, B 
                           => en, Y => n2276);
   U7220 : OAI2BB1X1 port map( A0N => n371, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_13_port, 
                           B0 => n2275, Y => n2293);
   U7221 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_12_port, B 
                           => en, Y => n2275);
   U7222 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_14_port, 
                           B0 => n2274, Y => n2292);
   U7223 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_13_port, B 
                           => en, Y => n2274);
   U7224 : OAI2BB1X1 port map( A0N => n372, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_15_port, 
                           B0 => n2273, Y => n2291);
   U7225 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_14_port, B 
                           => en, Y => n2273);
   U7226 : OAI2BB1X1 port map( A0N => n368, A1N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_16_port, 
                           B0 => n2272, Y => n2290);
   U7227 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_15_port, B 
                           => en, Y => n2272);
   U7228 : OAI2BB1X1 port map( A0N => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_17_port, 
                           A1N => n371, B0 => n2271, Y => n2289);
   U7229 : NAND2X1 port map( A => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_16_port, B 
                           => en, Y => n2271);
   U7230 : INVX1 port map( A => n3570, Y => n1451);
   U7231 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_11, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_11_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3570);
   U7232 : INVX1 port map( A => n3567, Y => n1447);
   U7233 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_8, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_8_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3567);
   U7234 : INVX1 port map( A => n3561, Y => n1441);
   U7235 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_2, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_2_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3561);
   U7236 : INVX1 port map( A => n3588, Y => n1432);
   U7237 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_11, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_11_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3588);
   U7238 : INVX1 port map( A => n3585, Y => n1428);
   U7239 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_8, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_8_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3585);
   U7240 : INVX1 port map( A => n3579, Y => n1422);
   U7241 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_2, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_2_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3579);
   U7242 : INVX1 port map( A => n3606, Y => n1413);
   U7243 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_11,
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_11_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3606);
   U7244 : INVX1 port map( A => n3603, Y => n1409);
   U7245 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_8, 
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_8_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3603);
   U7246 : INVX1 port map( A => n3597, Y => n1403);
   U7247 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_2, 
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_2_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3597);
   U7248 : INVX1 port map( A => n3624, Y => n1394);
   U7249 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_11,
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_11_port, 
                           B1 => n7, Y => n3624);
   U7250 : INVX1 port map( A => n3621, Y => n1390);
   U7251 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_8, 
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_8_port, 
                           B1 => n7, Y => n3621);
   U7252 : INVX1 port map( A => n3615, Y => n1384);
   U7253 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_2, 
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_2_port, 
                           B1 => n7, Y => n3615);
   U7254 : INVX1 port map( A => input_times_b0_div_componentxUDxn13, Y => n1275
                           );
   U7255 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_11, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_11_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn13);
   U7256 : INVX1 port map( A => input_times_b0_div_componentxUDxn10, Y => n1271
                           );
   U7257 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_8, A1 
                           => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_8_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn10);
   U7258 : INVX1 port map( A => input_times_b0_div_componentxUDxn4, Y => n1265)
                           ;
   U7259 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_2, A1 
                           => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_2_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn4);
   U7260 : INVX1 port map( A => n3576, Y => n1457);
   U7261 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_17, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_17_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3576);
   U7262 : INVX1 port map( A => n3575, Y => n1456);
   U7263 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_16, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_16_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3575);
   U7264 : INVX1 port map( A => n3573, Y => n1454);
   U7265 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_14, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_14_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3573);
   U7266 : INVX1 port map( A => n3572, Y => n1453);
   U7267 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_13, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_13_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3572);
   U7268 : INVX1 port map( A => n3571, Y => n1452);
   U7269 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_12, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_12_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3571);
   U7270 : INVX1 port map( A => n3569, Y => n1450);
   U7271 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_10, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_10_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3569);
   U7272 : INVX1 port map( A => n3566, Y => n1446);
   U7273 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_7, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_7_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3566);
   U7274 : INVX1 port map( A => n3564, Y => n1444);
   U7275 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_5, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_5_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3564);
   U7276 : INVX1 port map( A => n3563, Y => n1443);
   U7277 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_4, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_4_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3563);
   U7278 : INVX1 port map( A => n3562, Y => n1442);
   U7279 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_3, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_3_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3562);
   U7280 : INVX1 port map( A => n3560, Y => n1440);
   U7281 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_1, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_1_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3560);
   U7282 : INVX1 port map( A => n3559, Y => n1439);
   U7283 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_0_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3559);
   U7284 : INVX1 port map( A => n3594, Y => n1438);
   U7285 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_17, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_17_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3594);
   U7286 : INVX1 port map( A => n3593, Y => n1437);
   U7287 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_16, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_16_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3593);
   U7288 : INVX1 port map( A => n3591, Y => n1435);
   U7289 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_14, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_14_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3591);
   U7290 : INVX1 port map( A => n3590, Y => n1434);
   U7291 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_13, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_13_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3590);
   U7292 : INVX1 port map( A => n3589, Y => n1433);
   U7293 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_12, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_12_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3589);
   U7294 : INVX1 port map( A => n3587, Y => n1431);
   U7295 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_10, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_10_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3587);
   U7296 : INVX1 port map( A => n3584, Y => n1427);
   U7297 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_7, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_7_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3584);
   U7298 : INVX1 port map( A => n3582, Y => n1425);
   U7299 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_5, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_5_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3582);
   U7300 : INVX1 port map( A => n3581, Y => n1424);
   U7301 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_4, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_4_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3581);
   U7302 : INVX1 port map( A => n3580, Y => n1423);
   U7303 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_3, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_3_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3580);
   U7304 : INVX1 port map( A => n3578, Y => n1421);
   U7305 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_1, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_1_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3578);
   U7306 : INVX1 port map( A => n3577, Y => n1420);
   U7307 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_0_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3577);
   U7308 : INVX1 port map( A => n3612, Y => n1419);
   U7309 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_17,
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_17_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3612);
   U7310 : INVX1 port map( A => n3611, Y => n1418);
   U7311 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_16,
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_16_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3611);
   U7312 : INVX1 port map( A => n3609, Y => n1416);
   U7313 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_14,
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_14_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3609);
   U7314 : INVX1 port map( A => n3608, Y => n1415);
   U7315 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_13,
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_13_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3608);
   U7316 : INVX1 port map( A => n3607, Y => n1414);
   U7317 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_12,
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_12_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3607);
   U7318 : INVX1 port map( A => n3605, Y => n1412);
   U7319 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_10,
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_10_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3605);
   U7320 : INVX1 port map( A => n3602, Y => n1408);
   U7321 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_7, 
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_7_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3602);
   U7322 : INVX1 port map( A => n3600, Y => n1406);
   U7323 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_5, 
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_5_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3600);
   U7324 : INVX1 port map( A => n3599, Y => n1405);
   U7325 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_4, 
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_4_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3599);
   U7326 : INVX1 port map( A => n3598, Y => n1404);
   U7327 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_3, 
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_3_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3598);
   U7328 : INVX1 port map( A => n3596, Y => n1402);
   U7329 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_1, 
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_1_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3596);
   U7330 : INVX1 port map( A => n3595, Y => n1401);
   U7331 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_0_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3595);
   U7332 : INVX1 port map( A => n3630, Y => n1400);
   U7333 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_17,
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_17_port, 
                           B1 => n7, Y => n3630);
   U7334 : INVX1 port map( A => n3629, Y => n1399);
   U7335 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_16,
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_16_port, 
                           B1 => n7, Y => n3629);
   U7336 : INVX1 port map( A => n3627, Y => n1397);
   U7337 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_14,
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_14_port, 
                           B1 => n7, Y => n3627);
   U7338 : INVX1 port map( A => n3626, Y => n1396);
   U7339 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_13,
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_13_port, 
                           B1 => n7, Y => n3626);
   U7340 : INVX1 port map( A => n3625, Y => n1395);
   U7341 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_12,
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_12_port, 
                           B1 => n7, Y => n3625);
   U7342 : INVX1 port map( A => n3623, Y => n1393);
   U7343 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_10,
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_10_port, 
                           B1 => n7, Y => n3623);
   U7344 : INVX1 port map( A => n3620, Y => n1389);
   U7345 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_7, 
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_7_port, 
                           B1 => n7, Y => n3620);
   U7346 : INVX1 port map( A => n3618, Y => n1387);
   U7347 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_5, 
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_5_port, 
                           B1 => n7, Y => n3618);
   U7348 : INVX1 port map( A => n3617, Y => n1386);
   U7349 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_4, 
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_4_port, 
                           B1 => n7, Y => n3617);
   U7350 : INVX1 port map( A => n3616, Y => n1385);
   U7351 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_3, 
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_3_port, 
                           B1 => n7, Y => n3616);
   U7352 : INVX1 port map( A => n3614, Y => n1383);
   U7353 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_1, 
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_1_port, 
                           B1 => n7, Y => n3614);
   U7354 : INVX1 port map( A => n3613, Y => n1382);
   U7355 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_0_port, 
                           B1 => n7, Y => n3613);
   U7356 : INVX1 port map( A => input_times_b0_div_componentxUDxn19, Y => n1281
                           );
   U7357 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_17, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_17_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn19);
   U7358 : INVX1 port map( A => input_times_b0_div_componentxUDxn18, Y => n1280
                           );
   U7359 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_16, A1 
                           => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_16_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn18);
   U7360 : INVX1 port map( A => input_times_b0_div_componentxUDxn16, Y => n1278
                           );
   U7361 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_14, A1 
                           => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_14_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn16);
   U7362 : INVX1 port map( A => input_times_b0_div_componentxUDxn15, Y => n1277
                           );
   U7363 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_13, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_13_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn15);
   U7364 : INVX1 port map( A => input_times_b0_div_componentxUDxn14, Y => n1276
                           );
   U7365 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_12, A1 
                           => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_12_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn14);
   U7366 : INVX1 port map( A => input_times_b0_div_componentxUDxn12, Y => n1274
                           );
   U7367 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_10, A1 
                           => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_10_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn12);
   U7368 : INVX1 port map( A => input_times_b0_div_componentxUDxn9, Y => n1270)
                           ;
   U7369 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_7, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_7_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn9);
   U7370 : INVX1 port map( A => input_times_b0_div_componentxUDxn7, Y => n1268)
                           ;
   U7371 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_5, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_5_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn7);
   U7372 : INVX1 port map( A => input_times_b0_div_componentxUDxn6, Y => n1267)
                           ;
   U7373 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_4, A1 
                           => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_4_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn6);
   U7374 : INVX1 port map( A => input_times_b0_div_componentxUDxn5, Y => n1266)
                           ;
   U7375 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_3, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_3_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn5);
   U7376 : INVX1 port map( A => input_times_b0_div_componentxUDxn3, Y => n1264)
                           ;
   U7377 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_1, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_1_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn3);
   U7378 : INVX1 port map( A => input_times_b0_div_componentxUDxn1, Y => n1263)
                           ;
   U7379 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_inverted_0_port, 
                           A1 => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_0_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn1);
   U7380 : INVX1 port map( A => n3574, Y => n1455);
   U7381 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_15, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_15_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3574);
   U7382 : INVX1 port map( A => n3568, Y => n1449);
   U7383 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_9, 
                           A1 => n159, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_9_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3568);
   U7384 : INVX1 port map( A => n3565, Y => n1445);
   U7385 : AOI22X1 port map( A0 => 
                           input_p1_times_b1_div_componentxunsigned_output_6, 
                           A1 => n160, B0 => 
                           input_p1_times_b1_div_componentxUDxquotient_not_gated_6_port, 
                           B1 => 
                           input_p1_times_b1_div_componentxoutput_ready_signal,
                           Y => n3565);
   U7386 : INVX1 port map( A => n3592, Y => n1436);
   U7387 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_15, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_15_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3592);
   U7388 : INVX1 port map( A => n3586, Y => n1430);
   U7389 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_9, 
                           A1 => n157, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_9_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3586);
   U7390 : INVX1 port map( A => n3583, Y => n1426);
   U7391 : AOI22X1 port map( A0 => 
                           input_p2_times_b2_div_componentxunsigned_output_6, 
                           A1 => n158, B0 => 
                           input_p2_times_b2_div_componentxUDxquotient_not_gated_6_port, 
                           B1 => 
                           input_p2_times_b2_div_componentxoutput_ready_signal,
                           Y => n3583);
   U7392 : INVX1 port map( A => n3610, Y => n1417);
   U7393 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_15,
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_15_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3610);
   U7394 : INVX1 port map( A => n3604, Y => n1411);
   U7395 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_9, 
                           A1 => n155, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_9_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3604);
   U7396 : INVX1 port map( A => n3601, Y => n1407);
   U7397 : AOI22X1 port map( A0 => 
                           output_p1_times_a1_div_componentxunsigned_output_6, 
                           A1 => n156, B0 => 
                           output_p1_times_a1_div_componentxUDxquotient_not_gated_6_port, 
                           B1 => 
                           output_p1_times_a1_div_componentxoutput_ready_signal
                           , Y => n3601);
   U7398 : INVX1 port map( A => n3628, Y => n1398);
   U7399 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_15,
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_15_port, 
                           B1 => n7, Y => n3628);
   U7400 : INVX1 port map( A => n3622, Y => n1392);
   U7401 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_9, 
                           A1 => n153, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_9_port, 
                           B1 => n7, Y => n3622);
   U7402 : INVX1 port map( A => n3619, Y => n1388);
   U7403 : AOI22X1 port map( A0 => 
                           output_p2_times_a2_div_componentxunsigned_output_6, 
                           A1 => n154, B0 => 
                           output_p2_times_a2_div_componentxUDxquotient_not_gated_6_port, 
                           B1 => n7, Y => n3619);
   U7404 : INVX1 port map( A => input_times_b0_div_componentxUDxn17, Y => n1279
                           );
   U7405 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_15, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_15_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn17);
   U7406 : INVX1 port map( A => input_times_b0_div_componentxUDxn11, Y => n1273
                           );
   U7407 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_9, A1 
                           => n137, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_9_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn11);
   U7408 : INVX1 port map( A => input_times_b0_div_componentxUDxn8, Y => n1269)
                           ;
   U7409 : AOI22X1 port map( A0 => 
                           input_times_b0_div_componentxunsigned_output_6, A1 
                           => n138, B0 => 
                           input_times_b0_div_componentxUDxquotient_not_gated_6_port, 
                           B1 => n8, Y => input_times_b0_div_componentxUDxn8);
   U7410 : AOI22X1 port map( A0 => parameter_B0_div(2), A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_2_port
                           , B1 => n341, Y => input_times_b0_div_componentxn47)
                           ;
   U7411 : XNOR2X1 port map( A => parameter_B0_div(2), B => n3889, Y => 
                           input_times_b0_div_componentxinput_B_inverted_2_port
                           );
   U7412 : NOR2X1 port map( A => parameter_B0_div(0), B => parameter_B0_div(1),
                           Y => n3889);
   U7413 : AOI22X1 port map( A0 => parameter_B1_div(2), A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_2_port, 
                           B1 => n332, Y => n4225);
   U7414 : XNOR2X1 port map( A => parameter_B1_div(2), B => n3932, Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_2_port);
   U7415 : NOR2X1 port map( A => parameter_B1_div(0), B => parameter_B1_div(1),
                           Y => n3932);
   U7416 : AOI22X1 port map( A0 => parameter_B2_div(2), A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_2_port, 
                           B1 => n323, Y => n4281);
   U7417 : XNOR2X1 port map( A => parameter_B2_div(2), B => n3975, Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_2_port);
   U7418 : NOR2X1 port map( A => parameter_B2_div(0), B => parameter_B2_div(1),
                           Y => n3975);
   U7419 : AOI22X1 port map( A0 => parameter_A1_div(2), A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_2_port, 
                           B1 => n359, Y => n4335);
   U7420 : XNOR2X1 port map( A => parameter_A1_div(2), B => n4018, Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_2_port);
   U7421 : NOR2X1 port map( A => parameter_A1_div(0), B => parameter_A1_div(1),
                           Y => n4018);
   U7422 : AOI22X1 port map( A0 => parameter_A2_div(2), A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_2_port, 
                           B1 => n350, Y => n4391);
   U7423 : XNOR2X1 port map( A => parameter_A2_div(2), B => n4061, Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_2_port);
   U7424 : NOR2X1 port map( A => parameter_A2_div(0), B => parameter_A2_div(1),
                           Y => n4061);
   U7425 : AOI22X1 port map( A0 => parameter_B0_div(4), A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_4_port
                           , B1 => n341, Y => input_times_b0_div_componentxn49)
                           ;
   U7426 : XOR2X1 port map( A => n3887, B => parameter_B0_div(4), Y => 
                           input_times_b0_div_componentxinput_B_inverted_4_port
                           );
   U7427 : OR2X2 port map( A => parameter_B0_div(3), B => n3888, Y => n3887);
   U7428 : AOI22X1 port map( A0 => parameter_B1_div(4), A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_4_port, 
                           B1 => n332, Y => n4227);
   U7429 : XOR2X1 port map( A => n3930, B => parameter_B1_div(4), Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_4_port);
   U7430 : OR2X2 port map( A => parameter_B1_div(3), B => n3931, Y => n3930);
   U7431 : AOI22X1 port map( A0 => parameter_B2_div(4), A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_4_port, 
                           B1 => n323, Y => n4283);
   U7432 : XOR2X1 port map( A => n3973, B => parameter_B2_div(4), Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_4_port);
   U7433 : OR2X2 port map( A => parameter_B2_div(3), B => n3974, Y => n3973);
   U7434 : AOI22X1 port map( A0 => parameter_A1_div(4), A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_4_port, 
                           B1 => n359, Y => n4337);
   U7435 : XOR2X1 port map( A => n4016, B => parameter_A1_div(4), Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_4_port);
   U7436 : OR2X2 port map( A => parameter_A1_div(3), B => n4017, Y => n4016);
   U7437 : AOI22X1 port map( A0 => parameter_A2_div(4), A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_4_port, 
                           B1 => n350, Y => n4393);
   U7438 : XOR2X1 port map( A => n4059, B => parameter_A2_div(4), Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_4_port);
   U7439 : OR2X2 port map( A => parameter_A2_div(3), B => n4060, Y => n4059);
   U7440 : AOI22X1 port map( A0 => parameter_B0_div(6), A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_6_port
                           , B1 => n341, Y => input_times_b0_div_componentxn51)
                           ;
   U7441 : XOR2X1 port map( A => n3885, B => parameter_B0_div(6), Y => 
                           input_times_b0_div_componentxinput_B_inverted_6_port
                           );
   U7442 : OR2X2 port map( A => parameter_B0_div(5), B => n3886, Y => n3885);
   U7443 : AOI22X1 port map( A0 => parameter_B1_div(6), A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_6_port, 
                           B1 => n332, Y => n4229);
   U7444 : XOR2X1 port map( A => n3928, B => parameter_B1_div(6), Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_6_port);
   U7445 : OR2X2 port map( A => parameter_B1_div(5), B => n3929, Y => n3928);
   U7446 : AOI22X1 port map( A0 => parameter_B2_div(6), A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_6_port, 
                           B1 => n323, Y => n4285);
   U7447 : XOR2X1 port map( A => n3971, B => parameter_B2_div(6), Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_6_port);
   U7448 : OR2X2 port map( A => parameter_B2_div(5), B => n3972, Y => n3971);
   U7449 : AOI22X1 port map( A0 => parameter_A1_div(6), A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_6_port, 
                           B1 => n359, Y => n4339);
   U7450 : XOR2X1 port map( A => n4014, B => parameter_A1_div(6), Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_6_port);
   U7451 : OR2X2 port map( A => parameter_A1_div(5), B => n4015, Y => n4014);
   U7452 : AOI22X1 port map( A0 => parameter_A2_div(6), A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_6_port, 
                           B1 => n350, Y => n4395);
   U7453 : XOR2X1 port map( A => n4057, B => parameter_A2_div(6), Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_6_port);
   U7454 : OR2X2 port map( A => parameter_A2_div(5), B => n4058, Y => n4057);
   U7455 : AOI22X1 port map( A0 => parameter_B0_div(3), A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_3_port
                           , B1 => n341, Y => input_times_b0_div_componentxn48)
                           ;
   U7456 : XOR2X1 port map( A => n3888, B => parameter_B0_div(3), Y => 
                           input_times_b0_div_componentxinput_B_inverted_3_port
                           );
   U7457 : AOI22X1 port map( A0 => parameter_B1_div(3), A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_3_port, 
                           B1 => n332, Y => n4226);
   U7458 : XOR2X1 port map( A => n3931, B => parameter_B1_div(3), Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_3_port);
   U7459 : AOI22X1 port map( A0 => parameter_B2_div(3), A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_3_port, 
                           B1 => n323, Y => n4282);
   U7460 : XOR2X1 port map( A => n3974, B => parameter_B2_div(3), Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_3_port);
   U7461 : AOI22X1 port map( A0 => parameter_A1_div(3), A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_3_port, 
                           B1 => n359, Y => n4336);
   U7462 : XOR2X1 port map( A => n4017, B => parameter_A1_div(3), Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_3_port);
   U7463 : AOI22X1 port map( A0 => parameter_A2_div(3), A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_3_port, 
                           B1 => n350, Y => n4392);
   U7464 : XOR2X1 port map( A => n4060, B => parameter_A2_div(3), Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_3_port);
   U7465 : AOI22X1 port map( A0 => parameter_B0_div(5), A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_5_port
                           , B1 => n341, Y => input_times_b0_div_componentxn50)
                           ;
   U7466 : XOR2X1 port map( A => n3886, B => parameter_B0_div(5), Y => 
                           input_times_b0_div_componentxinput_B_inverted_5_port
                           );
   U7467 : AOI22X1 port map( A0 => parameter_B1_div(5), A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_5_port, 
                           B1 => n332, Y => n4228);
   U7468 : XOR2X1 port map( A => n3929, B => parameter_B1_div(5), Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_5_port);
   U7469 : AOI22X1 port map( A0 => parameter_B2_div(5), A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_5_port, 
                           B1 => n323, Y => n4284);
   U7470 : XOR2X1 port map( A => n3972, B => parameter_B2_div(5), Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_5_port);
   U7471 : AOI22X1 port map( A0 => parameter_A1_div(5), A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_5_port, 
                           B1 => n359, Y => n4338);
   U7472 : XOR2X1 port map( A => n4015, B => parameter_A1_div(5), Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_5_port);
   U7473 : AOI22X1 port map( A0 => parameter_A2_div(5), A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_5_port, 
                           B1 => n350, Y => n4394);
   U7474 : XOR2X1 port map( A => n4058, B => parameter_A2_div(5), Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_5_port);
   U7475 : INVX1 port map( A => input_times_b0_div_componentxn45, Y => n846);
   U7476 : AOI22X1 port map( A0 => parameter_B0_div(0), A1 => n342, B0 => 
                           parameter_B0_div(0), B1 => n341, Y => 
                           input_times_b0_div_componentxn45);
   U7477 : INVX1 port map( A => n4223, Y => n1005);
   U7478 : AOI22X1 port map( A0 => parameter_B1_div(0), A1 => n333, B0 => 
                           parameter_B1_div(0), B1 => n332, Y => n4223);
   U7479 : INVX1 port map( A => n4279, Y => n1164);
   U7480 : AOI22X1 port map( A0 => parameter_B2_div(0), A1 => n324, B0 => 
                           parameter_B2_div(0), B1 => n323, Y => n4279);
   U7481 : INVX1 port map( A => n4333, Y => n528);
   U7482 : AOI22X1 port map( A0 => parameter_A1_div(0), A1 => n360, B0 => 
                           parameter_A1_div(0), B1 => n359, Y => n4333);
   U7483 : INVX1 port map( A => n4389, Y => n687);
   U7484 : AOI22X1 port map( A0 => parameter_A2_div(0), A1 => n351, B0 => 
                           parameter_A2_div(0), B1 => n350, Y => n4389);
   U7485 : OR3XL port map( A => parameter_B1_mul(5), B => parameter_B1_mul(6), 
                           C => n3699, Y => n3697);
   U7486 : OR3XL port map( A => parameter_B2_mul(5), B => parameter_B2_mul(6), 
                           C => n3747, Y => n3745);
   U7487 : OR3XL port map( A => parameter_A2_mul(5), B => parameter_A2_mul(6), 
                           C => n3843, Y => n3841);
   U7488 : OR3XL port map( A => parameter_B0_mul(5), B => parameter_B0_mul(6), 
                           C => n3651, Y => n3649);
   U7489 : OR3XL port map( A => parameter_A1_mul(5), B => parameter_A1_mul(6), 
                           C => n3795, Y => n3793);
   U7490 : OR3XL port map( A => parameter_B0_div(5), B => parameter_B0_div(6), 
                           C => n3886, Y => n3884);
   U7491 : OR3XL port map( A => parameter_B1_div(5), B => parameter_B1_div(6), 
                           C => n3929, Y => n3927);
   U7492 : OR3XL port map( A => parameter_B2_div(5), B => parameter_B2_div(6), 
                           C => n3972, Y => n3970);
   U7493 : OR3XL port map( A => parameter_A1_div(5), B => parameter_A1_div(6), 
                           C => n4015, Y => n4013);
   U7494 : OR3XL port map( A => parameter_A2_div(5), B => parameter_A2_div(6), 
                           C => n4058, Y => n4056);
   U7495 : OR3XL port map( A => parameter_B1_mul(3), B => parameter_B1_mul(4), 
                           C => n3701, Y => n3699);
   U7496 : OR3XL port map( A => parameter_B2_mul(3), B => parameter_B2_mul(4), 
                           C => n3749, Y => n3747);
   U7497 : OR3XL port map( A => parameter_A2_mul(3), B => parameter_A2_mul(4), 
                           C => n3845, Y => n3843);
   U7498 : OR3XL port map( A => parameter_B0_mul(3), B => parameter_B0_mul(4), 
                           C => n3653, Y => n3651);
   U7499 : OR3XL port map( A => parameter_B0_div(3), B => parameter_B0_div(4), 
                           C => n3888, Y => n3886);
   U7500 : OR3XL port map( A => parameter_B1_div(3), B => parameter_B1_div(4), 
                           C => n3931, Y => n3929);
   U7501 : OR3XL port map( A => parameter_B2_div(3), B => parameter_B2_div(4), 
                           C => n3974, Y => n3972);
   U7502 : OR3XL port map( A => parameter_A1_mul(3), B => parameter_A1_mul(4), 
                           C => n3797, Y => n3795);
   U7503 : OR3XL port map( A => parameter_A1_div(3), B => parameter_A1_div(4), 
                           C => n4017, Y => n4015);
   U7504 : OR3XL port map( A => parameter_A2_div(3), B => parameter_A2_div(4), 
                           C => n4060, Y => n4058);
   U7505 : OR3XL port map( A => parameter_B1_mul(1), B => parameter_B1_mul(2), 
                           C => parameter_B1_mul(0), Y => n3701);
   U7506 : OR3XL port map( A => parameter_B2_mul(1), B => parameter_B2_mul(2), 
                           C => parameter_B2_mul(0), Y => n3749);
   U7507 : OR3XL port map( A => parameter_A1_mul(1), B => parameter_A1_mul(2), 
                           C => parameter_A1_mul(0), Y => n3797);
   U7508 : OR3XL port map( A => parameter_A2_mul(1), B => parameter_A2_mul(2), 
                           C => parameter_A2_mul(0), Y => n3845);
   U7509 : OR3XL port map( A => parameter_B0_mul(1), B => parameter_B0_mul(2), 
                           C => parameter_B0_mul(0), Y => n3653);
   U7510 : OR3XL port map( A => parameter_B0_div(1), B => parameter_B0_div(2), 
                           C => parameter_B0_div(0), Y => n3888);
   U7511 : OR3XL port map( A => parameter_B1_div(1), B => parameter_B1_div(2), 
                           C => parameter_B1_div(0), Y => n3931);
   U7512 : OR3XL port map( A => parameter_B2_div(1), B => parameter_B2_div(2), 
                           C => parameter_B2_div(0), Y => n3974);
   U7513 : OR3XL port map( A => parameter_A1_div(1), B => parameter_A1_div(2), 
                           C => parameter_A1_div(0), Y => n4017);
   U7514 : OR3XL port map( A => parameter_A2_div(1), B => parameter_A2_div(2), 
                           C => parameter_A2_div(0), Y => n4060);
   U7515 : BUFX3 port map( A => n4423, Y => n179);
   U7516 : AOI22X1 port map( A0 => parameter_B1_mul(0), A1 => n339, B0 => 
                           parameter_B1_mul(0), B1 => n336, Y => n4423);
   U7517 : BUFX3 port map( A => n4476, Y => n200);
   U7518 : AOI22X1 port map( A0 => parameter_B2_mul(0), A1 => n330, B0 => 
                           parameter_B2_mul(0), B1 => n327, Y => n4476);
   U7519 : BUFX3 port map( A => n4582, Y => n242);
   U7520 : AOI22X1 port map( A0 => parameter_A2_mul(0), A1 => n357, B0 => 
                           parameter_A2_mul(0), B1 => n354, Y => n4582);
   U7521 : BUFX3 port map( A => input_times_b0_mul_componentxn72, Y => n270);
   U7522 : AOI22X1 port map( A0 => parameter_B0_mul(0), A1 => n348, B0 => 
                           parameter_B0_mul(0), B1 => n345, Y => 
                           input_times_b0_mul_componentxn72);
   U7523 : BUFX3 port map( A => n4529, Y => n221);
   U7524 : AOI22X1 port map( A0 => parameter_A1_mul(0), A1 => n366, B0 => 
                           parameter_A1_mul(0), B1 => n363, Y => n4529);
   U7525 : BUFX3 port map( A => n4415, Y => n178);
   U7526 : AOI22X1 port map( A0 => parameter_B1_mul(1), A1 => n338, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_1_port, 
                           B1 => n335, Y => n4415);
   U7527 : XOR2X1 port map( A => parameter_B1_mul(1), B => parameter_B1_mul(0),
                           Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_1_port);
   U7528 : BUFX3 port map( A => n4468, Y => n199);
   U7529 : AOI22X1 port map( A0 => parameter_B2_mul(1), A1 => n329, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_1_port, 
                           B1 => n326, Y => n4468);
   U7530 : XOR2X1 port map( A => parameter_B2_mul(1), B => parameter_B2_mul(0),
                           Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_1_port);
   U7531 : BUFX3 port map( A => n4521, Y => n220);
   U7532 : AOI22X1 port map( A0 => parameter_A1_mul(1), A1 => n365, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_1_port, 
                           B1 => n362, Y => n4521);
   U7533 : XOR2X1 port map( A => parameter_A1_mul(1), B => parameter_A1_mul(0),
                           Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_1_port);
   U7534 : BUFX3 port map( A => n4574, Y => n241);
   U7535 : AOI22X1 port map( A0 => parameter_A2_mul(1), A1 => n356, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_1_port, 
                           B1 => n353, Y => n4574);
   U7536 : XOR2X1 port map( A => parameter_A2_mul(1), B => parameter_A2_mul(0),
                           Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_1_port);
   U7537 : BUFX3 port map( A => input_times_b0_mul_componentxn64, Y => n269);
   U7538 : AOI22X1 port map( A0 => parameter_B0_mul(1), A1 => n347, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_1_port
                           , B1 => n344, Y => input_times_b0_mul_componentxn64)
                           ;
   U7539 : XOR2X1 port map( A => parameter_B0_mul(1), B => parameter_B0_mul(0),
                           Y => 
                           input_times_b0_mul_componentxinput_B_inverted_1_port
                           );
   U7540 : BUFX3 port map( A => n4414, Y => n177);
   U7541 : AOI22X1 port map( A0 => parameter_B1_mul(2), A1 => n338, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_2_port, 
                           B1 => n335, Y => n4414);
   U7542 : XNOR2X1 port map( A => parameter_B1_mul(2), B => n3702, Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_2_port);
   U7543 : NOR2X1 port map( A => parameter_B1_mul(0), B => parameter_B1_mul(1),
                           Y => n3702);
   U7544 : BUFX3 port map( A => n4467, Y => n198);
   U7545 : AOI22X1 port map( A0 => parameter_B2_mul(2), A1 => n329, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_2_port, 
                           B1 => n326, Y => n4467);
   U7546 : XNOR2X1 port map( A => parameter_B2_mul(2), B => n3750, Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_2_port);
   U7547 : NOR2X1 port map( A => parameter_B2_mul(0), B => parameter_B2_mul(1),
                           Y => n3750);
   U7548 : BUFX3 port map( A => n4520, Y => n219);
   U7549 : AOI22X1 port map( A0 => parameter_A1_mul(2), A1 => n365, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_2_port, 
                           B1 => n362, Y => n4520);
   U7550 : XNOR2X1 port map( A => parameter_A1_mul(2), B => n3798, Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_2_port);
   U7551 : NOR2X1 port map( A => parameter_A1_mul(0), B => parameter_A1_mul(1),
                           Y => n3798);
   U7552 : BUFX3 port map( A => n4573, Y => n240);
   U7553 : AOI22X1 port map( A0 => parameter_A2_mul(2), A1 => n356, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_2_port, 
                           B1 => n353, Y => n4573);
   U7554 : XNOR2X1 port map( A => parameter_A2_mul(2), B => n3846, Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_2_port);
   U7555 : NOR2X1 port map( A => parameter_A2_mul(0), B => parameter_A2_mul(1),
                           Y => n3846);
   U7556 : BUFX3 port map( A => input_times_b0_mul_componentxn63, Y => n268);
   U7557 : AOI22X1 port map( A0 => parameter_B0_mul(2), A1 => n347, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_2_port
                           , B1 => n345, Y => input_times_b0_mul_componentxn63)
                           ;
   U7558 : XNOR2X1 port map( A => parameter_B0_mul(2), B => n3654, Y => 
                           input_times_b0_mul_componentxinput_B_inverted_2_port
                           );
   U7559 : NOR2X1 port map( A => parameter_B0_mul(0), B => parameter_B0_mul(1),
                           Y => n3654);
   U7560 : BUFX3 port map( A => n4413, Y => n176);
   U7561 : AOI22X1 port map( A0 => parameter_B1_mul(3), A1 => n339, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_3_port, 
                           B1 => n335, Y => n4413);
   U7562 : XOR2X1 port map( A => n3701, B => parameter_B1_mul(3), Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_3_port);
   U7563 : BUFX3 port map( A => n4466, Y => n197);
   U7564 : AOI22X1 port map( A0 => parameter_B2_mul(3), A1 => n330, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_3_port, 
                           B1 => n326, Y => n4466);
   U7565 : XOR2X1 port map( A => n3749, B => parameter_B2_mul(3), Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_3_port);
   U7566 : BUFX3 port map( A => n4519, Y => n218);
   U7567 : AOI22X1 port map( A0 => parameter_A1_mul(3), A1 => n366, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_3_port, 
                           B1 => n362, Y => n4519);
   U7568 : XOR2X1 port map( A => n3797, B => parameter_A1_mul(3), Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_3_port);
   U7569 : BUFX3 port map( A => n4572, Y => n239);
   U7570 : AOI22X1 port map( A0 => parameter_A2_mul(3), A1 => n357, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_3_port, 
                           B1 => n353, Y => n4572);
   U7571 : XOR2X1 port map( A => n3845, B => parameter_A2_mul(3), Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_3_port);
   U7572 : BUFX3 port map( A => input_times_b0_mul_componentxn62, Y => n267);
   U7573 : AOI22X1 port map( A0 => parameter_B0_mul(3), A1 => n348, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_3_port
                           , B1 => n344, Y => input_times_b0_mul_componentxn62)
                           ;
   U7574 : XOR2X1 port map( A => n3653, B => parameter_B0_mul(3), Y => 
                           input_times_b0_mul_componentxinput_B_inverted_3_port
                           );
   U7575 : INVX1 port map( A => en, Y => n368);
   U7576 : BUFX3 port map( A => n4412, Y => n175);
   U7577 : AOI22X1 port map( A0 => parameter_B1_mul(4), A1 => n338, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_4_port, 
                           B1 => n335, Y => n4412);
   U7578 : XOR2X1 port map( A => n3700, B => parameter_B1_mul(4), Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_4_port);
   U7579 : OR2X2 port map( A => parameter_B1_mul(3), B => n3701, Y => n3700);
   U7580 : BUFX3 port map( A => n4465, Y => n196);
   U7581 : AOI22X1 port map( A0 => parameter_B2_mul(4), A1 => n329, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_4_port, 
                           B1 => n326, Y => n4465);
   U7582 : XOR2X1 port map( A => n3748, B => parameter_B2_mul(4), Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_4_port);
   U7583 : OR2X2 port map( A => parameter_B2_mul(3), B => n3749, Y => n3748);
   U7584 : BUFX3 port map( A => n4518, Y => n217);
   U7585 : AOI22X1 port map( A0 => parameter_A1_mul(4), A1 => n365, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_4_port, 
                           B1 => n362, Y => n4518);
   U7586 : XOR2X1 port map( A => n3796, B => parameter_A1_mul(4), Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_4_port);
   U7587 : OR2X2 port map( A => parameter_A1_mul(3), B => n3797, Y => n3796);
   U7588 : BUFX3 port map( A => n4571, Y => n238);
   U7589 : AOI22X1 port map( A0 => parameter_A2_mul(4), A1 => n356, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_4_port, 
                           B1 => n353, Y => n4571);
   U7590 : XOR2X1 port map( A => n3844, B => parameter_A2_mul(4), Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_4_port);
   U7591 : OR2X2 port map( A => parameter_A2_mul(3), B => n3845, Y => n3844);
   U7592 : BUFX3 port map( A => input_times_b0_mul_componentxn61, Y => n266);
   U7593 : AOI22X1 port map( A0 => parameter_B0_mul(4), A1 => n347, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_4_port
                           , B1 => n344, Y => input_times_b0_mul_componentxn61)
                           ;
   U7594 : XOR2X1 port map( A => n3652, B => parameter_B0_mul(4), Y => 
                           input_times_b0_mul_componentxinput_B_inverted_4_port
                           );
   U7595 : OR2X2 port map( A => parameter_B0_mul(3), B => n3653, Y => n3652);
   U7596 : INVX1 port map( A => input_times_b0_div_componentxn46, Y => n847);
   U7597 : AOI22X1 port map( A0 => parameter_B0_div(1), A1 => n342, B0 => 
                           input_times_b0_div_componentxinput_B_inverted_1_port
                           , B1 => n341, Y => input_times_b0_div_componentxn46)
                           ;
   U7598 : XOR2X1 port map( A => parameter_B0_div(1), B => parameter_B0_div(0),
                           Y => 
                           input_times_b0_div_componentxinput_B_inverted_1_port
                           );
   U7599 : INVX1 port map( A => n4224, Y => n1006);
   U7600 : AOI22X1 port map( A0 => parameter_B1_div(1), A1 => n333, B0 => 
                           input_p1_times_b1_div_componentxinput_B_inverted_1_port, 
                           B1 => n332, Y => n4224);
   U7601 : XOR2X1 port map( A => parameter_B1_div(1), B => parameter_B1_div(0),
                           Y => 
                           input_p1_times_b1_div_componentxinput_B_inverted_1_port);
   U7602 : INVX1 port map( A => n4280, Y => n1165);
   U7603 : AOI22X1 port map( A0 => parameter_B2_div(1), A1 => n324, B0 => 
                           input_p2_times_b2_div_componentxinput_B_inverted_1_port, 
                           B1 => n323, Y => n4280);
   U7604 : XOR2X1 port map( A => parameter_B2_div(1), B => parameter_B2_div(0),
                           Y => 
                           input_p2_times_b2_div_componentxinput_B_inverted_1_port);
   U7605 : INVX1 port map( A => n4334, Y => n529);
   U7606 : AOI22X1 port map( A0 => parameter_A1_div(1), A1 => n360, B0 => 
                           output_p1_times_a1_div_componentxinput_B_inverted_1_port, 
                           B1 => n359, Y => n4334);
   U7607 : XOR2X1 port map( A => parameter_A1_div(1), B => parameter_A1_div(0),
                           Y => 
                           output_p1_times_a1_div_componentxinput_B_inverted_1_port);
   U7608 : INVX1 port map( A => n4390, Y => n688);
   U7609 : AOI22X1 port map( A0 => parameter_A2_div(1), A1 => n351, B0 => 
                           output_p2_times_a2_div_componentxinput_B_inverted_1_port, 
                           B1 => n350, Y => n4390);
   U7610 : XOR2X1 port map( A => parameter_A2_div(1), B => parameter_A2_div(0),
                           Y => 
                           output_p2_times_a2_div_componentxinput_B_inverted_1_port);
   U7611 : BUFX3 port map( A => n4411, Y => n174);
   U7612 : AOI22X1 port map( A0 => parameter_B1_mul(5), A1 => n339, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_5_port, 
                           B1 => n335, Y => n4411);
   U7613 : XOR2X1 port map( A => n3699, B => parameter_B1_mul(5), Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_5_port);
   U7614 : BUFX3 port map( A => n4464, Y => n195);
   U7615 : AOI22X1 port map( A0 => parameter_B2_mul(5), A1 => n330, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_5_port, 
                           B1 => n326, Y => n4464);
   U7616 : XOR2X1 port map( A => n3747, B => parameter_B2_mul(5), Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_5_port);
   U7617 : BUFX3 port map( A => n4517, Y => n216);
   U7618 : AOI22X1 port map( A0 => parameter_A1_mul(5), A1 => n366, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_5_port, 
                           B1 => n362, Y => n4517);
   U7619 : XOR2X1 port map( A => n3795, B => parameter_A1_mul(5), Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_5_port);
   U7620 : BUFX3 port map( A => n4570, Y => n237);
   U7621 : AOI22X1 port map( A0 => parameter_A2_mul(5), A1 => n357, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_5_port, 
                           B1 => n353, Y => n4570);
   U7622 : XOR2X1 port map( A => n3843, B => parameter_A2_mul(5), Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_5_port);
   U7623 : BUFX3 port map( A => input_times_b0_mul_componentxn60, Y => n265);
   U7624 : AOI22X1 port map( A0 => parameter_B0_mul(5), A1 => n348, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_5_port
                           , B1 => n344, Y => input_times_b0_mul_componentxn60)
                           ;
   U7625 : XOR2X1 port map( A => n3651, B => parameter_B0_mul(5), Y => 
                           input_times_b0_mul_componentxinput_B_inverted_5_port
                           );
   U7626 : INVX1 port map( A => n337, Y => n336);
   U7627 : INVX1 port map( A => n328, Y => n327);
   U7628 : INVX1 port map( A => n355, Y => n354);
   U7629 : INVX1 port map( A => n346, Y => n345);
   U7630 : INVX1 port map( A => n364, Y => n363);
   U7631 : BUFX3 port map( A => n4410, Y => n173);
   U7632 : AOI22X1 port map( A0 => parameter_B1_mul(6), A1 => n338, B0 => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_6_port, 
                           B1 => n335, Y => n4410);
   U7633 : XOR2X1 port map( A => n3698, B => parameter_B1_mul(6), Y => 
                           input_p1_times_b1_mul_componentxinput_B_inverted_6_port);
   U7634 : OR2X2 port map( A => parameter_B1_mul(5), B => n3699, Y => n3698);
   U7635 : BUFX3 port map( A => n4463, Y => n194);
   U7636 : AOI22X1 port map( A0 => parameter_B2_mul(6), A1 => n329, B0 => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_6_port, 
                           B1 => n326, Y => n4463);
   U7637 : XOR2X1 port map( A => n3746, B => parameter_B2_mul(6), Y => 
                           input_p2_times_b2_mul_componentxinput_B_inverted_6_port);
   U7638 : OR2X2 port map( A => parameter_B2_mul(5), B => n3747, Y => n3746);
   U7639 : BUFX3 port map( A => n4516, Y => n215);
   U7640 : AOI22X1 port map( A0 => parameter_A1_mul(6), A1 => n365, B0 => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_6_port, 
                           B1 => n362, Y => n4516);
   U7641 : XOR2X1 port map( A => n3794, B => parameter_A1_mul(6), Y => 
                           output_p1_times_a1_mul_componentxinput_B_inverted_6_port);
   U7642 : OR2X2 port map( A => parameter_A1_mul(5), B => n3795, Y => n3794);
   U7643 : BUFX3 port map( A => n4569, Y => n236);
   U7644 : AOI22X1 port map( A0 => parameter_A2_mul(6), A1 => n356, B0 => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_6_port, 
                           B1 => n353, Y => n4569);
   U7645 : XOR2X1 port map( A => n3842, B => parameter_A2_mul(6), Y => 
                           output_p2_times_a2_mul_componentxinput_B_inverted_6_port);
   U7646 : OR2X2 port map( A => parameter_A2_mul(5), B => n3843, Y => n3842);
   U7647 : BUFX3 port map( A => input_times_b0_mul_componentxn59, Y => n264);
   U7648 : AOI22X1 port map( A0 => parameter_B0_mul(6), A1 => n347, B0 => 
                           input_times_b0_mul_componentxinput_B_inverted_6_port
                           , B1 => n344, Y => input_times_b0_mul_componentxn59)
                           ;
   U7649 : XOR2X1 port map( A => n3650, B => parameter_B0_mul(6), Y => 
                           input_times_b0_mul_componentxinput_B_inverted_6_port
                           );
   U7650 : OR2X2 port map( A => parameter_B0_mul(5), B => n3651, Y => n3650);
   U7651 : INVX1 port map( A => input_signal(7), Y => n1174);
   U7652 : INVX1 port map( A => parameter_B0_div(7), Y => n342);
   U7653 : INVX1 port map( A => parameter_B1_div(7), Y => n333);
   U7654 : INVX1 port map( A => parameter_B2_div(7), Y => n324);
   U7655 : INVX1 port map( A => parameter_A1_div(7), Y => n360);
   U7656 : INVX1 port map( A => parameter_A2_div(7), Y => n351);
   U7657 : INVX1 port map( A => parameter_B1_mul(7), Y => n339);
   U7658 : INVX1 port map( A => parameter_B2_mul(7), Y => n330);
   U7659 : INVX1 port map( A => parameter_A2_mul(7), Y => n357);
   U7660 : INVX1 port map( A => parameter_A1_mul(7), Y => n366);
   U7661 : INVX1 port map( A => parameter_B0_mul(7), Y => n348);
   U7662 : INVX1 port map( A => parameter_B1_mul(7), Y => n337);
   U7663 : INVX1 port map( A => parameter_B2_mul(7), Y => n328);
   U7664 : INVX1 port map( A => parameter_A2_mul(7), Y => n355);
   U7665 : INVX1 port map( A => parameter_B0_mul(7), Y => n346);
   U7666 : INVX1 port map( A => parameter_A1_mul(7), Y => n364);
   U7667 : INVX1 port map( A => parameter_B1_mul(7), Y => n338);
   U7668 : INVX1 port map( A => parameter_B2_mul(7), Y => n329);
   U7669 : INVX1 port map( A => parameter_A1_mul(7), Y => n365);
   U7670 : INVX1 port map( A => parameter_A2_mul(7), Y => n356);
   U7671 : INVX1 port map( A => parameter_B0_mul(7), Y => n347);

end SYN_flow_arch;
